
module datapath ( clock, reset, inputSRAM_Data, graphRead1_DataInput, 
        graphRead2_DataInput, workRead1_DataInput, workRead2_DataInput, 
        inputSRAM_Addr, graphRead1_Addr, graphRead2_Addr, workWrite_Dist, 
        workWrite_Pred, workRead1_Addr, workRead2_Addr, workWrite_Addr, 
        work_WE, outputWrite_Data, outputWrite_Addr, output_WE, state, 
        graphData1_Zero_reg, iterDone, iterStop, negCycle, zeroFlag, 
        outputWriteDone, goS8 );
  input [7:0] inputSRAM_Data;
  input [127:0] graphRead1_DataInput;
  input [127:0] graphRead2_DataInput;
  input [127:0] workRead1_DataInput;
  input [127:0] workRead2_DataInput;
  output [9:0] inputSRAM_Addr;
  output [12:0] graphRead1_Addr;
  output [12:0] graphRead2_Addr;
  output [16:0] workWrite_Dist;
  output [7:0] workWrite_Pred;
  output [12:0] workRead1_Addr;
  output [12:0] workRead2_Addr;
  output [12:0] workWrite_Addr;
  output [15:0] outputWrite_Data;
  output [13:0] outputWrite_Addr;
  input [4:0] state;
  input clock, reset;
  output work_WE, output_WE, graphData1_Zero_reg, iterDone, iterStop, negCycle,
         zeroFlag, outputWriteDone, goS8;
  wire   U3_U3_DATA6_1, U3_U3_DATA6_2, U3_U3_DATA6_3, U3_U3_DATA6_4,
         U3_U3_DATA6_5, U3_U3_DATA6_6, U3_U3_DATA6_7, U3_U3_DATA6_8,
         U3_U3_DATA6_9, U3_U3_DATA6_10, U3_U6_Z_0, U3_U6_DATA4_1,
         U3_U6_DATA4_5, U3_U6_DATA4_6, U3_U6_DATA4_7, U113_DATA2_0,
         U113_DATA2_1, U113_DATA2_2, U113_DATA2_3, U113_DATA2_4, U113_DATA2_5,
         U113_DATA2_6, U113_DATA2_7, U112_DATA1_0, U112_DATA1_1, U112_DATA1_2,
         U112_DATA1_3, U112_DATA1_4, U112_DATA1_5, U112_DATA1_6, U112_DATA1_7,
         U112_DATA1_8, U112_DATA1_9, U112_DATA1_10, U112_DATA1_11,
         U112_DATA1_12, U112_DATA1_13, U112_DATA1_14, U112_DATA1_15,
         U112_DATA1_16, U97_DATA4_0, U97_DATA4_1, U97_DATA4_2, U97_DATA4_3,
         U97_DATA4_4, U97_DATA4_5, U97_DATA4_6, U97_DATA4_7, U97_DATA3_3,
         U97_DATA3_4, U97_DATA3_5, U97_DATA3_6, U97_DATA3_7, U97_DATA2_0,
         U97_DATA2_1, U97_DATA2_2, U97_DATA2_3, U97_DATA2_4, U97_DATA2_5,
         U97_DATA2_6, U97_DATA2_7, U92_DATA2_0, U92_DATA2_1, U92_DATA2_2,
         U92_DATA2_3, U92_DATA2_4, U92_DATA2_5, U92_DATA2_6, U92_DATA2_7,
         U91_DATA2_0, U91_DATA2_1, U91_DATA2_2, U91_DATA2_3, U91_DATA2_4,
         U91_DATA2_5, U91_DATA2_6, U91_DATA2_7, U38_DATA6_0, U38_DATA6_1,
         U38_DATA6_2, U38_DATA6_3, U38_DATA6_4, U38_DATA6_5, U38_DATA6_6,
         U38_DATA6_7, U38_DATA5_0, U38_DATA5_1, U38_DATA5_2, U38_DATA5_3,
         U38_DATA5_4, U38_DATA5_5, U38_DATA5_6, U38_DATA5_7, U38_DATA4_0,
         U38_DATA4_1, U38_DATA4_2, U38_DATA4_3, U38_DATA4_4, U38_DATA4_5,
         U38_DATA4_6, U38_DATA4_7, U38_DATA3_0, U38_DATA3_1, U38_DATA3_2,
         U38_DATA3_3, U38_DATA3_4, U38_DATA3_5, U38_DATA3_6, U38_DATA3_7,
         U38_DATA2_0, U38_DATA2_1, U38_DATA2_2, U38_DATA2_3, U38_DATA2_4,
         U38_DATA2_5, U38_DATA2_6, U38_DATA2_7, U38_DATA1_0, U38_DATA1_1,
         U38_DATA1_2, U38_DATA1_3, U38_DATA1_4, U38_DATA1_5, U38_DATA1_6,
         U38_DATA1_7, U37_DATA6_0, U37_DATA6_1, U37_DATA6_2, U37_DATA6_3,
         U37_DATA6_4, U37_DATA6_5, U37_DATA6_6, U37_DATA6_7, U37_DATA5_0,
         U37_DATA5_1, U37_DATA5_2, U37_DATA5_3, U37_DATA5_4, U37_DATA5_5,
         U37_DATA5_6, U37_DATA5_7, U37_DATA2_0, U37_DATA2_1, U37_DATA2_2,
         U37_DATA2_3, U37_DATA2_4, U37_DATA2_5, U37_DATA2_6, U37_DATA2_7,
         U37_DATA1_0, U37_DATA1_1, U37_DATA1_2, U37_DATA1_3, U37_DATA1_4,
         U37_DATA1_5, U37_DATA1_6, U37_DATA1_7, U16_DATA2_1, U16_DATA2_2,
         U16_DATA2_3, U16_DATA2_4, U16_DATA2_5, U16_DATA2_6, U16_DATA2_7,
         U16_DATA2_8, U16_DATA2_9, U16_DATA2_10, U16_DATA2_11, U16_DATA2_12,
         U16_DATA2_13, U8_DATA3_1, U8_DATA3_2, U8_DATA3_3, U8_DATA3_4,
         U8_DATA3_5, U8_DATA3_6, U8_DATA3_7, sub_387_carry_2_,
         sub_387_carry_3_, sub_387_carry_4_, sub_387_carry_5_,
         sub_387_carry_6_, sub_387_carry_7_, sub_387_A_0_, sub_387_A_1_,
         sub_387_A_2_, sub_387_A_3_, sub_387_A_4_, sub_387_A_5_, sub_387_A_6_,
         sub_387_A_7_, r572_A_0_, r572_A_1_, r572_A_2_, eq_565_B_7_,
         eq_565_B_6_, eq_565_B_5_, eq_565_B_4_, eq_565_B_3_, eq_565_B_2_,
         eq_565_B_1_, eq_565_B_0_, mult_add_378_aco_a_2_,
         mult_add_378_aco_a_1_, mult_add_378_aco_a_0_, add_118_A_16_, n2, n3,
         n4, n5, n6, n7, n8, n9, n11, n13, n15, n17, n19, n21, n23, n25, n27,
         n29, n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n125, n127, n129, n131, n133, n135, n137, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n273, n275,
         n277, n279, n281, n283, n285, n287, n289, n291, n293, n294, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n391, n392,
         n393, n394, n395, n396, n397, n398, n416, n417, n418, n421, n424,
         n425, n430, n431, n432, n433, n434, n438, n439, n440, n441, n442,
         n443, n444, n445, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n563, n564, n575, n577, n578, n579, n594,
         n595, n600, n606, n612, n618, n624, n630, n637, n682, n725, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n828, n830, n831, n832, n834, n835, n836, n837,
         n842, n844, n845, n849, n893, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n981, n982, n983, n988, n989, n991, n993, n995,
         n997, n999, n1001, n1003, n1005, n1006, n1011, n1013, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1025, n1026, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1040, n1041, n1042, n1047,
         n1049, n1050, n1051, n1054, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, net10760, net10761, net10766, net10803, net10805,
         net10828, net10830, net10834, net10835, net10839, net10840, net10842,
         net10844, net10849, net10850, net10863, net10867, net10881, net10884,
         net10885, net10887, net10893, net10899, net10903, net10907, net10911,
         net10915, net10919, net10923, net10927, net10931, net10939, net10940,
         net10942, net10943, net10950, net11085, net11093, net11113, net11117,
         net11119, net11121, net11126, net11131, net11136, net11164, net11165,
         net11170, net11171, net11175, net11186, net11226, net11227, net11236,
         net11292, net11309, net11311, net11312, net11316, net11334, net11335,
         net11368, net11375, net11384, net11387, net11399, net11403, net11417,
         net11425, net11431, net11450, net11454, net11458, net11466, net11498,
         net11516, net11518, net11520, net11581, net11584, net11586, net11590,
         net11592, net11605, net11609, net11623, net11631, net11632, net11636,
         net11640, net11644, net11648, net11682, net11670, net11668, net11700,
         net11696, net11694, net11742, net11750, net11754, net11856, net11894,
         net12569, net12566, net12578, net12590, net12597, net12622, net12620,
         net12639, net12649, net12722, net12724, net12730, net12766, net12921,
         net12938, net12936, net12943, net12959, net12968, net12979, net13012,
         net13011, net13034, net13039, net13049, net13082, net11195, net11162,
         n669, n668, n667, n666, n665, n664, n663, n662, net11474, net11473,
         net11405, net11475, net10765, net15569, net17911, net17910, net10841,
         net10837, n251, net17864, net10913, net10898, net10846, net10937,
         net10930, net10922, net10921, net10920, net10941, net10936, net10851,
         net10847, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160;
  wire   [11:2] r520_carry;

  HA_X1 r520_U1_1_1 ( .A(graphRead1_Addr[1]), .B(graphRead1_Addr[0]), .CO(
        r520_carry[2]), .S(U3_U3_DATA6_1) );
  HA_X1 r520_U1_1_2 ( .A(graphRead1_Addr[2]), .B(r520_carry[2]), .CO(
        r520_carry[3]), .S(U3_U3_DATA6_2) );
  HA_X1 r520_U1_1_3 ( .A(graphRead1_Addr[3]), .B(r520_carry[3]), .CO(
        r520_carry[4]), .S(U3_U3_DATA6_3) );
  HA_X1 r520_U1_1_4 ( .A(graphRead1_Addr[4]), .B(r520_carry[4]), .CO(
        r520_carry[5]), .S(U3_U3_DATA6_4) );
  HA_X1 r520_U1_1_5 ( .A(graphRead1_Addr[5]), .B(r520_carry[5]), .CO(
        r520_carry[6]), .S(U3_U3_DATA6_5) );
  HA_X1 r520_U1_1_6 ( .A(graphRead1_Addr[6]), .B(r520_carry[6]), .CO(
        r520_carry[7]), .S(U3_U3_DATA6_6) );
  HA_X1 r520_U1_1_7 ( .A(graphRead1_Addr[7]), .B(r520_carry[7]), .CO(
        r520_carry[8]), .S(U3_U3_DATA6_7) );
  HA_X1 r520_U1_1_8 ( .A(graphRead1_Addr[8]), .B(r520_carry[8]), .CO(
        r520_carry[9]), .S(U3_U3_DATA6_8) );
  HA_X1 r520_U1_1_9 ( .A(graphRead1_Addr[9]), .B(r520_carry[9]), .CO(
        r520_carry[10]), .S(U3_U3_DATA6_9) );
  HA_X1 r520_U1_1_10 ( .A(graphRead1_Addr[10]), .B(r520_carry[10]), .CO(
        r520_carry[11]), .S(U3_U3_DATA6_10) );
  XNOR2_X2 sub_387_U1_A_1 ( .A(sub_387_A_1_), .B(sub_387_A_0_), .ZN(U8_DATA3_1) );
  XNOR2_X2 sub_387_U1_A_2 ( .A(sub_387_A_2_), .B(sub_387_carry_2_), .ZN(
        U8_DATA3_2) );
  OR2_X1 sub_387_U1_B_2 ( .A1(sub_387_A_2_), .A2(sub_387_carry_2_), .ZN(
        sub_387_carry_3_) );
  XNOR2_X2 sub_387_U1_A_3 ( .A(sub_387_A_3_), .B(sub_387_carry_3_), .ZN(
        U8_DATA3_3) );
  OR2_X1 sub_387_U1_B_3 ( .A1(sub_387_A_3_), .A2(sub_387_carry_3_), .ZN(
        sub_387_carry_4_) );
  XNOR2_X2 sub_387_U1_A_4 ( .A(sub_387_A_4_), .B(sub_387_carry_4_), .ZN(
        U8_DATA3_4) );
  OR2_X1 sub_387_U1_B_4 ( .A1(sub_387_A_4_), .A2(sub_387_carry_4_), .ZN(
        sub_387_carry_5_) );
  XNOR2_X2 sub_387_U1_A_5 ( .A(sub_387_A_5_), .B(sub_387_carry_5_), .ZN(
        U8_DATA3_5) );
  OR2_X1 sub_387_U1_B_5 ( .A1(sub_387_A_5_), .A2(sub_387_carry_5_), .ZN(
        sub_387_carry_6_) );
  XNOR2_X2 sub_387_U1_A_6 ( .A(sub_387_A_6_), .B(sub_387_carry_6_), .ZN(
        U8_DATA3_6) );
  OR2_X1 sub_387_U1_B_6 ( .A1(sub_387_A_6_), .A2(sub_387_carry_6_), .ZN(
        sub_387_carry_7_) );
  XNOR2_X2 sub_387_U1_A_7 ( .A(sub_387_A_7_), .B(sub_387_carry_7_), .ZN(
        U8_DATA3_7) );
  DFF_X2 daughterCount_reg_0_ ( .D(n1404), .CK(clock), .Q(net12938), .QN(n337)
         );
  DFF_X2 inputSRAM_Addr_reg_1_ ( .D(n1395), .CK(clock), .Q(inputSRAM_Addr[1]), 
        .QN(n268) );
  DFF_X2 inputSRAM_Addr_reg_2_ ( .D(n1394), .CK(clock), .Q(inputSRAM_Addr[2]), 
        .QN(n266) );
  DFF_X2 inputSRAM_Addr_reg_3_ ( .D(n1393), .CK(clock), .Q(inputSRAM_Addr[3]), 
        .QN(n264) );
  DFF_X2 inputSRAM_Addr_reg_4_ ( .D(n1392), .CK(clock), .Q(inputSRAM_Addr[4]), 
        .QN(n262) );
  DFF_X2 inputSRAM_Addr_reg_5_ ( .D(n1391), .CK(clock), .Q(inputSRAM_Addr[5]), 
        .QN(n260) );
  DFF_X2 inputSRAM_Addr_reg_6_ ( .D(n1390), .CK(clock), .Q(inputSRAM_Addr[6]), 
        .QN(n258) );
  DFF_X2 inputSRAM_Addr_reg_7_ ( .D(n1389), .CK(clock), .Q(inputSRAM_Addr[7]), 
        .QN(n256) );
  DFF_X2 totalVertex_reg_1_ ( .D(n1341), .CK(clock), .QN(n86) );
  DFF_X2 graphRead1_Addr_reg_8_ ( .D(n1326), .CK(clock), .Q(graphRead1_Addr[8]), .QN(n277) );
  DFF_X2 graphRead1_Addr_reg_9_ ( .D(n1325), .CK(clock), .Q(graphRead1_Addr[9]), .QN(n275) );
  DFF_X2 graphRead1_Addr_reg_10_ ( .D(n1324), .CK(clock), .Q(
        graphRead1_Addr[10]), .QN(n273) );
  DFF_X2 graphRead1_Addr_reg_11_ ( .D(n1323), .CK(clock), .Q(
        graphRead1_Addr[11]), .QN(n271) );
  DFF_X2 graphRead1_Addr_reg_12_ ( .D(n1322), .CK(clock), .Q(
        graphRead1_Addr[12]), .QN(n270) );
  DFF_X2 totalVertex_reg_0_ ( .D(n1342), .CK(clock), .QN(n87) );
  DFF_X2 vertexCount_reg_1_ ( .D(n1333), .CK(clock), .Q(sub_387_A_1_), .QN(n41) );
  DFF_X2 vertexCount_reg_2_ ( .D(n1332), .CK(clock), .Q(sub_387_A_2_), .QN(n40) );
  DFF_X2 vertexCount_reg_5_ ( .D(n1329), .CK(clock), .Q(sub_387_A_5_), .QN(n37) );
  DFF_X2 vertexCount_reg_6_ ( .D(n1328), .CK(clock), .Q(sub_387_A_6_), .QN(n36) );
  DFF_X2 vertexCount_reg_7_ ( .D(n1327), .CK(clock), .Q(sub_387_A_7_), .QN(n35) );
  DFF_X2 inputSRAM_Addr_reg_8_ ( .D(n1388), .CK(clock), .Q(inputSRAM_Addr[8]), 
        .QN(n254) );
  DFF_X2 inputSRAM_Addr_reg_9_ ( .D(n1387), .CK(clock), .Q(inputSRAM_Addr[9]), 
        .QN(n252) );
  DFF_X2 inputSRAM_Addr_reg_0_ ( .D(n1396), .CK(clock), .Q(inputSRAM_Addr[0]), 
        .QN(n269) );
  DFF_X2 workRead1_Dist_reg_16_ ( .D(n1320), .CK(clock), .Q(add_118_A_16_), 
        .QN(n2478) );
  DFF_X2 outputWrite_Data_reg_15_ ( .D(n1288), .CK(clock), .Q(
        outputWrite_Data[15]), .QN(n366) );
  DFF_X2 workRead1_Dist_reg_14_ ( .D(n1318), .CK(clock), .Q(U91_DATA2_6) );
  DFF_X2 outputWrite_Data_reg_14_ ( .D(n1289), .CK(clock), .Q(
        outputWrite_Data[14]), .QN(n367) );
  DFF_X2 outputWrite_Data_reg_13_ ( .D(n1290), .CK(clock), .Q(
        outputWrite_Data[13]), .QN(n368) );
  DFF_X2 outputWrite_Data_reg_12_ ( .D(n1291), .CK(clock), .Q(
        outputWrite_Data[12]), .QN(n369) );
  DFF_X2 outputWrite_Data_reg_11_ ( .D(n1292), .CK(clock), .Q(
        outputWrite_Data[11]), .QN(n370) );
  DFF_X2 outputWrite_Data_reg_10_ ( .D(n1293), .CK(clock), .Q(
        outputWrite_Data[10]), .QN(n371) );
  DFF_X2 outputWrite_Data_reg_9_ ( .D(n1294), .CK(clock), .Q(
        outputWrite_Data[9]), .QN(n372) );
  DFF_X2 outputWrite_Data_reg_8_ ( .D(n1295), .CK(clock), .Q(
        outputWrite_Data[8]), .QN(n373) );
  DFF_X2 workRead1_Dist_reg_7_ ( .D(n1311), .CK(clock), .Q(U92_DATA2_7), .QN(
        n2475) );
  DFF_X2 outputWrite_Data_reg_7_ ( .D(n1296), .CK(clock), .Q(
        outputWrite_Data[7]), .QN(n374) );
  DFF_X2 outputWrite_Data_reg_6_ ( .D(n1297), .CK(clock), .Q(
        outputWrite_Data[6]), .QN(n375) );
  DFF_X2 outputWrite_Data_reg_5_ ( .D(n1298), .CK(clock), .Q(
        outputWrite_Data[5]), .QN(n376) );
  DFF_X2 outputWrite_Data_reg_4_ ( .D(n1299), .CK(clock), .Q(
        outputWrite_Data[4]), .QN(n377) );
  DFF_X2 workRead1_Dist_reg_3_ ( .D(n1307), .CK(clock), .Q(U92_DATA2_3), .QN(
        n2476) );
  DFF_X2 outputWrite_Data_reg_3_ ( .D(n1300), .CK(clock), .Q(
        outputWrite_Data[3]), .QN(n378) );
  DFF_X2 workRead1_Dist_reg_2_ ( .D(n1306), .CK(clock), .Q(U92_DATA2_2), .QN(
        n2487) );
  DFF_X2 outputWrite_Data_reg_2_ ( .D(n1301), .CK(clock), .Q(
        outputWrite_Data[2]), .QN(n379) );
  DFF_X2 workRead1_Dist_reg_1_ ( .D(n1305), .CK(clock), .Q(U92_DATA2_1), .QN(
        n2496) );
  DFF_X2 outputWrite_Data_reg_1_ ( .D(n1302), .CK(clock), .Q(
        outputWrite_Data[1]), .QN(n380) );
  DFF_X2 workRead1_Dist_reg_0_ ( .D(n1304), .CK(clock), .Q(U92_DATA2_0) );
  DFF_X2 outputWrite_Data_reg_0_ ( .D(n1303), .CK(clock), .Q(
        outputWrite_Data[0]), .QN(n381) );
  DFF_X2 vertexAddress_reg_1_ ( .D(n1270), .CK(clock), .Q(graphRead2_Addr[1]), 
        .QN(n349) );
  DFF_X2 iterationCount_reg_1_ ( .D(n1283), .CK(clock), .QN(n33) );
  DFF_X2 vertexAddress_reg_2_ ( .D(n1269), .CK(clock), .Q(graphRead2_Addr[2]), 
        .QN(n348) );
  DFF_X2 iterationCount_reg_2_ ( .D(n1282), .CK(clock), .QN(n31) );
  DFF_X2 vertexAddress_reg_3_ ( .D(n1268), .CK(clock), .Q(graphRead2_Addr[3]), 
        .QN(n347) );
  DFF_X2 iterationCount_reg_3_ ( .D(n1281), .CK(clock), .QN(n29) );
  DFF_X2 vertexAddress_reg_4_ ( .D(n1267), .CK(clock), .Q(graphRead2_Addr[4]), 
        .QN(n346) );
  DFF_X2 iterationCount_reg_4_ ( .D(n1280), .CK(clock), .QN(n27) );
  DFF_X2 vertexAddress_reg_5_ ( .D(n1266), .CK(clock), .Q(graphRead2_Addr[5]), 
        .QN(n345) );
  DFF_X2 iterationCount_reg_5_ ( .D(n1279), .CK(clock), .QN(n25) );
  DFF_X2 vertexAddress_reg_6_ ( .D(n1265), .CK(clock), .Q(graphRead2_Addr[6]), 
        .QN(n344) );
  DFF_X2 iterationCount_reg_6_ ( .D(n1278), .CK(clock), .QN(n23) );
  DFF_X2 vertexAddress_reg_7_ ( .D(n1264), .CK(clock), .Q(graphRead2_Addr[7]), 
        .QN(n343) );
  DFF_X2 iterationCount_reg_7_ ( .D(n1277), .CK(clock), .QN(n21) );
  DFF_X2 vertexAddress_reg_8_ ( .D(n1263), .CK(clock), .Q(graphRead2_Addr[8]), 
        .QN(n342) );
  DFF_X2 iterationCount_reg_8_ ( .D(n1276), .CK(clock), .QN(n19) );
  DFF_X2 vertexAddress_reg_9_ ( .D(n1262), .CK(clock), .Q(graphRead2_Addr[9]), 
        .QN(n341) );
  DFF_X2 iterationCount_reg_9_ ( .D(n1275), .CK(clock), .QN(n17) );
  DFF_X2 vertexAddress_reg_10_ ( .D(n1261), .CK(clock), .Q(graphRead2_Addr[10]), .QN(n340) );
  DFF_X2 iterationCount_reg_10_ ( .D(n1274), .CK(clock), .QN(n15) );
  DFF_X2 vertexAddress_reg_11_ ( .D(n1260), .CK(clock), .Q(graphRead2_Addr[11]), .QN(n339) );
  DFF_X2 iterationCount_reg_11_ ( .D(n1273), .CK(clock), .QN(n13) );
  DFF_X2 vertexAddress_reg_12_ ( .D(n1259), .CK(clock), .Q(graphRead2_Addr[12]), .QN(n338) );
  DFF_X2 iterationCount_reg_12_ ( .D(n1272), .CK(clock), .QN(n11) );
  DFF_X2 vertexAddress_reg_0_ ( .D(n1271), .CK(clock), .Q(graphRead2_Addr[0]), 
        .QN(n350) );
  DFF_X2 iterationCount_reg_0_ ( .D(n1284), .CK(clock), .Q(n2641), .QN(n34) );
  DFF_X2 workRead2_Addr_reg_3_ ( .D(n1159), .CK(clock), .Q(workRead2_Addr[3]), 
        .QN(n100) );
  DFF_X2 workRead2_Addr_reg_4_ ( .D(n1158), .CK(clock), .Q(workRead2_Addr[4]), 
        .QN(n99) );
  DFF_X2 workRead2_Addr_reg_5_ ( .D(n1157), .CK(clock), .Q(workRead2_Addr[5]), 
        .QN(n98) );
  DFF_X2 workRead2_Addr_reg_6_ ( .D(n1156), .CK(clock), .Q(workRead2_Addr[6]), 
        .QN(n97) );
  DFF_X2 workRead2_Addr_reg_7_ ( .D(n1155), .CK(clock), .Q(workRead2_Addr[7]), 
        .QN(n96) );
  DFF_X2 workRead2_Addr_reg_0_ ( .D(n1162), .CK(clock), .Q(workRead2_Addr[0]), 
        .QN(n103) );
  DFF_X2 workRead2_Addr_reg_1_ ( .D(n1161), .CK(clock), .Q(workRead2_Addr[1]), 
        .QN(n102) );
  DFF_X2 workRead2_Addr_reg_2_ ( .D(n1160), .CK(clock), .Q(workRead2_Addr[2]), 
        .QN(n101) );
  NAND2_X2 U20 ( .A1(workWrite_Addr[7]), .A2(n3157), .ZN(n579) );
  NAND2_X2 U27 ( .A1(workWrite_Addr[6]), .A2(n3157), .ZN(n595) );
  NOR3_X2 U178 ( .A1(n727), .A2(n728), .A3(n729), .ZN(n725) );
  OAI22_X2 U179 ( .A1(n187), .A2(n730), .B1(n203), .B2(n731), .ZN(n729) );
  OAI22_X2 U180 ( .A1(n219), .A2(n732), .B1(n235), .B2(n733), .ZN(n728) );
  OAI221_X2 U181 ( .B1(n139), .B2(n734), .C1(n104), .C2(n735), .A(n736), .ZN(
        n727) );
  NOR3_X2 U184 ( .A1(n739), .A2(n740), .A3(n741), .ZN(n738) );
  OAI22_X2 U185 ( .A1(n188), .A2(n730), .B1(n204), .B2(n731), .ZN(n741) );
  OAI22_X2 U186 ( .A1(n220), .A2(n732), .B1(n236), .B2(n733), .ZN(n740) );
  OAI221_X2 U187 ( .B1(n140), .B2(n734), .C1(n105), .C2(n735), .A(n742), .ZN(
        n739) );
  NOR3_X2 U190 ( .A1(n744), .A2(n745), .A3(n746), .ZN(n743) );
  OAI22_X2 U191 ( .A1(n189), .A2(n730), .B1(n205), .B2(n731), .ZN(n746) );
  OAI22_X2 U192 ( .A1(n221), .A2(n732), .B1(n237), .B2(n733), .ZN(n745) );
  OAI221_X2 U193 ( .B1(n141), .B2(n734), .C1(n106), .C2(n735), .A(n747), .ZN(
        n744) );
  NOR3_X2 U196 ( .A1(n749), .A2(n750), .A3(n751), .ZN(n748) );
  OAI22_X2 U197 ( .A1(n190), .A2(n730), .B1(n206), .B2(n731), .ZN(n751) );
  OAI22_X2 U198 ( .A1(n222), .A2(n732), .B1(n238), .B2(n733), .ZN(n750) );
  OAI221_X2 U199 ( .B1(n142), .B2(n734), .C1(n107), .C2(n735), .A(n752), .ZN(
        n749) );
  NOR3_X2 U202 ( .A1(n754), .A2(n755), .A3(n756), .ZN(n753) );
  OAI22_X2 U203 ( .A1(n191), .A2(n730), .B1(n207), .B2(n731), .ZN(n756) );
  OAI22_X2 U204 ( .A1(n223), .A2(n732), .B1(n239), .B2(n733), .ZN(n755) );
  OAI221_X2 U205 ( .B1(n143), .B2(n734), .C1(n108), .C2(n735), .A(n757), .ZN(
        n754) );
  NOR3_X2 U208 ( .A1(n759), .A2(n760), .A3(n761), .ZN(n758) );
  OAI22_X2 U209 ( .A1(n192), .A2(n730), .B1(n208), .B2(n731), .ZN(n761) );
  OAI22_X2 U210 ( .A1(n224), .A2(n732), .B1(n240), .B2(n733), .ZN(n760) );
  OAI221_X2 U211 ( .B1(n144), .B2(n734), .C1(n109), .C2(n735), .A(n762), .ZN(
        n759) );
  NOR3_X2 U214 ( .A1(n764), .A2(n765), .A3(n766), .ZN(n763) );
  OAI22_X2 U215 ( .A1(n193), .A2(n730), .B1(n209), .B2(n731), .ZN(n766) );
  OAI22_X2 U216 ( .A1(n225), .A2(n732), .B1(n241), .B2(n733), .ZN(n765) );
  OAI221_X2 U217 ( .B1(n145), .B2(n734), .C1(n110), .C2(n735), .A(n767), .ZN(
        n764) );
  NOR3_X2 U221 ( .A1(n769), .A2(n770), .A3(n771), .ZN(n768) );
  OAI22_X2 U222 ( .A1(n194), .A2(n730), .B1(n210), .B2(n731), .ZN(n771) );
  NAND3_X2 U223 ( .A1(r572_A_0_), .A2(n60), .A3(r572_A_2_), .ZN(n731) );
  NAND3_X2 U224 ( .A1(n61), .A2(n60), .A3(r572_A_2_), .ZN(n730) );
  OAI22_X2 U225 ( .A1(n226), .A2(n732), .B1(n242), .B2(n733), .ZN(n770) );
  NAND2_X2 U226 ( .A1(r572_A_2_), .A2(n772), .ZN(n733) );
  NAND3_X2 U227 ( .A1(r572_A_1_), .A2(n61), .A3(r572_A_2_), .ZN(n732) );
  OAI221_X2 U228 ( .B1(n146), .B2(n734), .C1(n111), .C2(n735), .A(n773), .ZN(
        n769) );
  NOR3_X2 U230 ( .A1(r572_A_0_), .A2(r572_A_2_), .A3(n60), .ZN(n737) );
  NAND3_X2 U231 ( .A1(n60), .A2(n59), .A3(r572_A_0_), .ZN(n734) );
  OAI221_X2 U402 ( .B1(n2494), .B2(n830), .C1(n424), .C2(n366), .A(n831), .ZN(
        n1288) );
  OAI221_X2 U403 ( .B1(n2556), .B2(n830), .C1(n424), .C2(n367), .A(n831), .ZN(
        n1289) );
  OAI221_X2 U404 ( .B1(n2497), .B2(n830), .C1(n424), .C2(n368), .A(n831), .ZN(
        n1290) );
  OAI221_X2 U405 ( .B1(n2492), .B2(n830), .C1(n424), .C2(n369), .A(n831), .ZN(
        n1291) );
  OAI221_X2 U406 ( .B1(n2495), .B2(n830), .C1(n424), .C2(n370), .A(n831), .ZN(
        n1292) );
  OAI221_X2 U407 ( .B1(n2491), .B2(n830), .C1(n424), .C2(n371), .A(n831), .ZN(
        n1293) );
  OAI221_X2 U408 ( .B1(n2474), .B2(n830), .C1(n424), .C2(n372), .A(n831), .ZN(
        n1294) );
  OAI221_X2 U409 ( .B1(n2498), .B2(n830), .C1(n424), .C2(n373), .A(n831), .ZN(
        n1295) );
  OAI221_X2 U410 ( .B1(n2475), .B2(n830), .C1(n424), .C2(n374), .A(n832), .ZN(
        n1296) );
  AOI221_X2 U411 ( .B1(U97_DATA3_7), .B2(n3158), .C1(U97_DATA4_7), .C2(n834), 
        .A(n70), .ZN(n832) );
  OAI221_X2 U412 ( .B1(n2493), .B2(n830), .C1(n424), .C2(n375), .A(n835), .ZN(
        n1297) );
  AOI221_X2 U413 ( .B1(U97_DATA3_6), .B2(n3158), .C1(U97_DATA4_6), .C2(n834), 
        .A(n70), .ZN(n835) );
  OAI221_X2 U414 ( .B1(n2481), .B2(n830), .C1(n424), .C2(n376), .A(n836), .ZN(
        n1298) );
  AOI221_X2 U415 ( .B1(U97_DATA3_5), .B2(n3158), .C1(U97_DATA4_5), .C2(n834), 
        .A(n70), .ZN(n836) );
  OAI221_X2 U416 ( .B1(n2490), .B2(n830), .C1(n424), .C2(n377), .A(n837), .ZN(
        n1299) );
  AOI221_X2 U417 ( .B1(U97_DATA3_4), .B2(n3158), .C1(U97_DATA4_4), .C2(n834), 
        .A(n70), .ZN(n837) );
  NOR2_X2 U427 ( .A1(zeroFlag), .A2(n844), .ZN(n842) );
  NOR2_X2 U428 ( .A1(n845), .A2(net11648), .ZN(n834) );
  OAI22_X2 U503 ( .A1(n425), .A2(n365), .B1(outputWrite_Addr[0]), .B2(n907), 
        .ZN(n1321) );
  NOR4_X2 U506 ( .A1(n912), .A2(outputWrite_Addr[3]), .A3(outputWrite_Addr[5]), 
        .A4(outputWrite_Addr[4]), .ZN(n911) );
  NOR4_X2 U507 ( .A1(n913), .A2(outputWrite_Addr[0]), .A3(outputWrite_Addr[11]), .A4(outputWrite_Addr[10]), .ZN(n910) );
  NAND4_X2 U544 ( .A1(n937), .A2(n938), .A3(n939), .A4(n940), .ZN(n936) );
  NOR4_X2 U545 ( .A1(graphRead1_DataInput[125]), .A2(graphRead1_DataInput[124]), .A3(graphRead1_DataInput[123]), .A4(graphRead1_DataInput[122]), .ZN(n940) );
  NOR4_X2 U546 ( .A1(graphRead1_DataInput[121]), .A2(graphRead1_DataInput[120]), .A3(graphRead1_DataInput[119]), .A4(graphRead1_DataInput[118]), .ZN(n939) );
  NOR4_X2 U547 ( .A1(graphRead1_DataInput[117]), .A2(graphRead1_DataInput[116]), .A3(graphRead1_DataInput[115]), .A4(graphRead1_DataInput[114]), .ZN(n938) );
  NOR4_X2 U548 ( .A1(graphRead1_DataInput[113]), .A2(graphRead1_DataInput[112]), .A3(graphRead1_DataInput[111]), .A4(graphRead1_DataInput[110]), .ZN(n937) );
  NAND4_X2 U549 ( .A1(n941), .A2(n942), .A3(n943), .A4(n944), .ZN(n935) );
  NOR4_X2 U550 ( .A1(graphRead1_DataInput[26]), .A2(graphRead1_DataInput[25]), 
        .A3(graphRead1_DataInput[24]), .A4(graphRead1_DataInput[23]), .ZN(n944) );
  NOR4_X2 U551 ( .A1(graphRead1_DataInput[22]), .A2(graphRead1_DataInput[21]), 
        .A3(graphRead1_DataInput[20]), .A4(graphRead1_DataInput[19]), .ZN(n943) );
  NOR4_X2 U552 ( .A1(graphRead1_DataInput[18]), .A2(graphRead1_DataInput[17]), 
        .A3(graphRead1_DataInput[16]), .A4(graphRead1_DataInput[15]), .ZN(n942) );
  NOR4_X2 U553 ( .A1(graphRead1_DataInput[14]), .A2(graphRead1_DataInput[13]), 
        .A3(graphRead1_DataInput[127]), .A4(graphRead1_DataInput[126]), .ZN(
        n941) );
  NAND4_X2 U554 ( .A1(n945), .A2(n946), .A3(n947), .A4(n948), .ZN(n934) );
  NOR4_X2 U555 ( .A1(graphRead1_DataInput[65]), .A2(graphRead1_DataInput[64]), 
        .A3(graphRead1_DataInput[9]), .A4(graphRead1_DataInput[8]), .ZN(n948)
         );
  NOR4_X2 U556 ( .A1(graphRead1_DataInput[7]), .A2(graphRead1_DataInput[6]), 
        .A3(graphRead1_DataInput[5]), .A4(graphRead1_DataInput[4]), .ZN(n947)
         );
  NOR4_X2 U557 ( .A1(graphRead1_DataInput[3]), .A2(graphRead1_DataInput[2]), 
        .A3(graphRead1_DataInput[12]), .A4(graphRead1_DataInput[11]), .ZN(n946) );
  NOR4_X2 U558 ( .A1(graphRead1_DataInput[10]), .A2(graphRead1_DataInput[1]), 
        .A3(graphRead1_DataInput[0]), .A4(n637), .ZN(n945) );
  NAND4_X2 U559 ( .A1(n949), .A2(n950), .A3(n951), .A4(n952), .ZN(n933) );
  NOR4_X2 U560 ( .A1(graphRead1_DataInput[109]), .A2(graphRead1_DataInput[108]), .A3(graphRead1_DataInput[107]), .A4(graphRead1_DataInput[106]), .ZN(n952) );
  NOR4_X2 U561 ( .A1(graphRead1_DataInput[105]), .A2(graphRead1_DataInput[104]), .A3(graphRead1_DataInput[103]), .A4(graphRead1_DataInput[102]), .ZN(n951) );
  NOR4_X2 U562 ( .A1(graphRead1_DataInput[101]), .A2(graphRead1_DataInput[100]), .A3(graphRead1_DataInput[71]), .A4(graphRead1_DataInput[70]), .ZN(n950) );
  NOR4_X2 U563 ( .A1(graphRead1_DataInput[69]), .A2(graphRead1_DataInput[68]), 
        .A3(graphRead1_DataInput[67]), .A4(graphRead1_DataInput[66]), .ZN(n949) );
  NAND4_X2 U564 ( .A1(n957), .A2(n958), .A3(n959), .A4(n960), .ZN(n956) );
  NOR4_X2 U565 ( .A1(graphRead1_DataInput[82]), .A2(graphRead1_DataInput[81]), 
        .A3(graphRead1_DataInput[80]), .A4(graphRead1_DataInput[79]), .ZN(n960) );
  NOR4_X2 U566 ( .A1(graphRead1_DataInput[78]), .A2(graphRead1_DataInput[77]), 
        .A3(graphRead1_DataInput[76]), .A4(graphRead1_DataInput[75]), .ZN(n959) );
  NOR4_X2 U567 ( .A1(graphRead1_DataInput[74]), .A2(graphRead1_DataInput[73]), 
        .A3(graphRead1_DataInput[72]), .A4(graphRead1_DataInput[63]), .ZN(n958) );
  NOR4_X2 U568 ( .A1(graphRead1_DataInput[62]), .A2(graphRead1_DataInput[61]), 
        .A3(graphRead1_DataInput[60]), .A4(graphRead1_DataInput[59]), .ZN(n957) );
  NAND4_X2 U569 ( .A1(n961), .A2(n962), .A3(n963), .A4(n964), .ZN(n955) );
  NOR4_X2 U570 ( .A1(n965), .A2(graphRead1_DataInput[97]), .A3(
        graphRead1_DataInput[99]), .A4(graphRead1_DataInput[98]), .ZN(n964) );
  NOR4_X2 U571 ( .A1(graphRead1_DataInput[94]), .A2(graphRead1_DataInput[93]), 
        .A3(graphRead1_DataInput[92]), .A4(graphRead1_DataInput[91]), .ZN(n963) );
  NOR4_X2 U572 ( .A1(graphRead1_DataInput[90]), .A2(graphRead1_DataInput[89]), 
        .A3(graphRead1_DataInput[88]), .A4(graphRead1_DataInput[87]), .ZN(n962) );
  NOR4_X2 U573 ( .A1(graphRead1_DataInput[86]), .A2(graphRead1_DataInput[85]), 
        .A3(graphRead1_DataInput[84]), .A4(graphRead1_DataInput[83]), .ZN(n961) );
  NAND4_X2 U574 ( .A1(n966), .A2(n967), .A3(n968), .A4(n969), .ZN(n954) );
  NOR4_X2 U575 ( .A1(graphRead1_DataInput[42]), .A2(graphRead1_DataInput[41]), 
        .A3(graphRead1_DataInput[40]), .A4(graphRead1_DataInput[39]), .ZN(n969) );
  NOR4_X2 U576 ( .A1(graphRead1_DataInput[38]), .A2(graphRead1_DataInput[37]), 
        .A3(graphRead1_DataInput[36]), .A4(graphRead1_DataInput[35]), .ZN(n968) );
  NOR4_X2 U577 ( .A1(graphRead1_DataInput[34]), .A2(graphRead1_DataInput[33]), 
        .A3(graphRead1_DataInput[32]), .A4(graphRead1_DataInput[31]), .ZN(n967) );
  NOR4_X2 U578 ( .A1(graphRead1_DataInput[30]), .A2(graphRead1_DataInput[29]), 
        .A3(graphRead1_DataInput[28]), .A4(graphRead1_DataInput[27]), .ZN(n966) );
  NAND4_X2 U579 ( .A1(n970), .A2(n971), .A3(n972), .A4(n973), .ZN(n953) );
  NOR4_X2 U580 ( .A1(graphRead1_DataInput[58]), .A2(graphRead1_DataInput[57]), 
        .A3(graphRead1_DataInput[56]), .A4(graphRead1_DataInput[55]), .ZN(n973) );
  NOR4_X2 U581 ( .A1(graphRead1_DataInput[54]), .A2(graphRead1_DataInput[53]), 
        .A3(graphRead1_DataInput[52]), .A4(graphRead1_DataInput[51]), .ZN(n972) );
  NOR4_X2 U582 ( .A1(graphRead1_DataInput[50]), .A2(graphRead1_DataInput[49]), 
        .A3(graphRead1_DataInput[48]), .A4(graphRead1_DataInput[47]), .ZN(n971) );
  NOR4_X2 U583 ( .A1(graphRead1_DataInput[46]), .A2(graphRead1_DataInput[45]), 
        .A3(graphRead1_DataInput[44]), .A4(graphRead1_DataInput[43]), .ZN(n970) );
  NOR2_X2 U597 ( .A1(n337), .A2(n336), .ZN(n983) );
  NAND2_X2 U625 ( .A1(workRead1_Addr[0]), .A2(n991), .ZN(n1006) );
  NAND2_X2 U626 ( .A1(reset), .A2(n54), .ZN(n989) );
  NAND3_X2 U650 ( .A1(n982), .A2(n337), .A3(U3_U6_DATA4_1), .ZN(n981) );
  NAND2_X2 U655 ( .A1(n772), .A2(n59), .ZN(n774) );
  NOR2_X2 U656 ( .A1(n60), .A2(n61), .ZN(n772) );
  NAND2_X2 U658 ( .A1(n1020), .A2(n1021), .ZN(n1019) );
  NOR2_X2 U659 ( .A1(n55), .A2(n1018), .ZN(n1017) );
  NOR2_X2 U660 ( .A1(n59), .A2(n1022), .ZN(n1018) );
  XNOR2_X2 U663 ( .A(n60), .B(r572_A_0_), .ZN(n1025) );
  NOR2_X2 U666 ( .A1(n55), .A2(n1021), .ZN(n1026) );
  NOR2_X2 U667 ( .A1(n60), .A2(n1022), .ZN(n1021) );
  NOR2_X2 U670 ( .A1(n61), .A2(n1022), .ZN(n1020) );
  NAND2_X2 U673 ( .A1(workRead1_DataInput[0]), .A2(n849), .ZN(n1029) );
  NAND2_X2 U675 ( .A1(workRead1_DataInput[1]), .A2(n849), .ZN(n1030) );
  NAND2_X2 U677 ( .A1(workRead1_DataInput[2]), .A2(n849), .ZN(n1031) );
  NAND2_X2 U679 ( .A1(workRead1_DataInput[3]), .A2(n849), .ZN(n1032) );
  NAND2_X2 U681 ( .A1(workRead1_DataInput[4]), .A2(n849), .ZN(n1033) );
  NAND2_X2 U683 ( .A1(workRead1_DataInput[5]), .A2(n849), .ZN(n1034) );
  NAND2_X2 U685 ( .A1(workRead1_DataInput[6]), .A2(n849), .ZN(n1035) );
  NAND2_X2 U687 ( .A1(workRead1_DataInput[7]), .A2(n849), .ZN(n1036) );
  OAI22_X2 U693 ( .A1(n1041), .A2(n254), .B1(n1042), .B2(n253), .ZN(n1388) );
  OAI22_X2 U694 ( .A1(n1041), .A2(n256), .B1(n1042), .B2(n255), .ZN(n1389) );
  OAI22_X2 U695 ( .A1(n1041), .A2(n258), .B1(n1042), .B2(n257), .ZN(n1390) );
  OAI22_X2 U696 ( .A1(n1041), .A2(n260), .B1(n1042), .B2(n259), .ZN(n1391) );
  OAI22_X2 U697 ( .A1(n1041), .A2(n262), .B1(n1042), .B2(n261), .ZN(n1392) );
  OAI22_X2 U698 ( .A1(n1041), .A2(n264), .B1(n1042), .B2(n263), .ZN(n1393) );
  OAI22_X2 U699 ( .A1(n1041), .A2(n266), .B1(n1042), .B2(n265), .ZN(n1394) );
  OAI22_X2 U700 ( .A1(n1041), .A2(n268), .B1(n1042), .B2(n267), .ZN(n1395) );
  OAI22_X2 U701 ( .A1(n1041), .A2(n269), .B1(U3_U6_Z_0), .B2(n1042), .ZN(n1396) );
  OAI22_X2 U717 ( .A1(n1047), .A2(n95), .B1(n1049), .B2(n3090), .ZN(n1405) );
  OAI22_X2 U718 ( .A1(n1047), .A2(n94), .B1(n1049), .B2(n3089), .ZN(n1406) );
  OAI22_X2 U719 ( .A1(n1047), .A2(n93), .B1(n1049), .B2(n3088), .ZN(n1407) );
  OAI22_X2 U720 ( .A1(n1047), .A2(n92), .B1(n1049), .B2(n434), .ZN(n1408) );
  OAI22_X2 U721 ( .A1(n1047), .A2(n91), .B1(n1049), .B2(n433), .ZN(n1409) );
  OAI22_X2 U722 ( .A1(n1047), .A2(n90), .B1(n1049), .B2(n432), .ZN(n1410) );
  OAI22_X2 U723 ( .A1(n1047), .A2(n89), .B1(n1049), .B2(n431), .ZN(n1411) );
  OAI22_X2 U724 ( .A1(n1047), .A2(n88), .B1(n1049), .B2(n430), .ZN(n1412) );
  NAND2_X2 U725 ( .A1(reset), .A2(n1047), .ZN(n1049) );
  NAND2_X2 U726 ( .A1(n1050), .A2(n1051), .ZN(n1413) );
  OAI22_X2 U737 ( .A1(n3098), .A2(n1058), .B1(n3090), .B2(n1059), .ZN(n1414)
         );
  OAI22_X2 U738 ( .A1(n3100), .A2(n1058), .B1(n3089), .B2(n1059), .ZN(n1415)
         );
  OAI22_X2 U739 ( .A1(n3102), .A2(n1058), .B1(n3088), .B2(n1059), .ZN(n1416)
         );
  OAI22_X2 U740 ( .A1(n3104), .A2(n1058), .B1(n434), .B2(n1059), .ZN(n1417) );
  OAI22_X2 U741 ( .A1(n3106), .A2(n1058), .B1(n433), .B2(n1059), .ZN(n1418) );
  OAI22_X2 U742 ( .A1(n3108), .A2(n1058), .B1(n432), .B2(n1059), .ZN(n1419) );
  OAI22_X2 U743 ( .A1(n3110), .A2(n1058), .B1(n431), .B2(n1059), .ZN(n1420) );
  OAI22_X2 U744 ( .A1(n3112), .A2(n1058), .B1(n430), .B2(n1059), .ZN(n1421) );
  NAND2_X2 U745 ( .A1(reset), .A2(n1058), .ZN(n1059) );
  NAND4_X2 U749 ( .A1(n434), .A2(n433), .A3(n1064), .A4(n432), .ZN(n1062) );
  NOR2_X2 U750 ( .A1(inputSRAM_Data[7]), .A2(inputSRAM_Data[6]), .ZN(n1064) );
  NOR4_X2 U751 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(negCycle)
         );
  NAND3_X2 U753 ( .A1(n27), .A2(n25), .A3(n29), .ZN(n1066) );
  NAND4_X2 U754 ( .A1(n23), .A2(n21), .A3(n19), .A4(n17), .ZN(n1065) );
  NOR4_X2 U755 ( .A1(n1069), .A2(n1070), .A3(sub_387_A_4_), .A4(sub_387_A_3_), 
        .ZN(iterDone) );
  NAND3_X2 U756 ( .A1(n36), .A2(n35), .A3(n37), .ZN(n1070) );
  NAND4_X2 U757 ( .A1(sub_387_A_0_), .A2(n828), .A3(n41), .A4(n40), .ZN(n1069)
         );
  NOR4_X2 U758 ( .A1(U97_DATA2_7), .A2(U97_DATA2_6), .A3(U97_DATA2_5), .A4(
        U97_DATA2_4), .ZN(n1072) );
  NOR4_X2 U759 ( .A1(U97_DATA2_3), .A2(U97_DATA2_2), .A3(U97_DATA2_1), .A4(
        U97_DATA2_0), .ZN(n1071) );
  NOR2_X2 U761 ( .A1(n337), .A2(n1073), .ZN(n828) );
  NOR2_X2 U762 ( .A1(n1074), .A2(n1075), .ZN(outputWriteDone) );
  NAND4_X2 U763 ( .A1(n1076), .A2(n1077), .A3(n1078), .A4(n1079), .ZN(n1075)
         );
  XNOR2_X2 U764 ( .A(eq_565_B_4_), .B(U97_DATA4_4), .ZN(n1079) );
  XNOR2_X2 U765 ( .A(eq_565_B_5_), .B(U97_DATA4_5), .ZN(n1078) );
  XNOR2_X2 U766 ( .A(eq_565_B_6_), .B(U97_DATA4_6), .ZN(n1077) );
  XNOR2_X2 U767 ( .A(eq_565_B_7_), .B(U97_DATA4_7), .ZN(n1076) );
  NAND4_X2 U768 ( .A1(n1080), .A2(n1081), .A3(n1082), .A4(n1083), .ZN(n1074)
         );
  XNOR2_X2 U769 ( .A(eq_565_B_0_), .B(U97_DATA4_0), .ZN(n1083) );
  XNOR2_X2 U770 ( .A(eq_565_B_1_), .B(U97_DATA4_1), .ZN(n1082) );
  XNOR2_X2 U771 ( .A(eq_565_B_2_), .B(U97_DATA4_2), .ZN(n1081) );
  XNOR2_X2 U772 ( .A(eq_565_B_3_), .B(U97_DATA4_3), .ZN(n1080) );
  AND3_X2 U776 ( .A1(n1054), .A2(n575), .A3(state[4]), .ZN(n1057) );
  NOR2_X2 U788 ( .A1(net11644), .A2(state[3]), .ZN(n1011) );
  NAND2_X2 U871 ( .A1(n982), .A2(n336), .ZN(n1073) );
  AND4_X2 U872 ( .A1(n334), .A2(n333), .A3(n335), .A4(n1120), .ZN(n982) );
  NOR3_X2 U873 ( .A1(U3_U6_DATA4_5), .A2(U3_U6_DATA4_7), .A3(U3_U6_DATA4_6), 
        .ZN(n1120) );
  INV_X4 U895 ( .A(n1019), .ZN(n57) );
  INV_X4 U896 ( .A(n774), .ZN(n58) );
  INV_X4 U898 ( .A(n1060), .ZN(n71) );
  INV_X4 U1006 ( .A(n893), .ZN(n351) );
  INV_X4 U1007 ( .A(n906), .ZN(n352) );
  INV_X4 U1008 ( .A(n905), .ZN(n353) );
  INV_X4 U1009 ( .A(n904), .ZN(n354) );
  INV_X4 U1010 ( .A(n903), .ZN(n355) );
  INV_X4 U1011 ( .A(n902), .ZN(n356) );
  INV_X4 U1012 ( .A(n901), .ZN(n357) );
  INV_X4 U1013 ( .A(n900), .ZN(n358) );
  INV_X4 U1014 ( .A(n899), .ZN(n359) );
  INV_X4 U1015 ( .A(n898), .ZN(n360) );
  INV_X4 U1016 ( .A(n897), .ZN(n361) );
  INV_X4 U1017 ( .A(n896), .ZN(n362) );
  INV_X4 U1018 ( .A(n895), .ZN(n363) );
  INV_X4 U1022 ( .A(n1061), .ZN(n421) );
  INV_X4 U1031 ( .A(inputSRAM_Data[7]), .ZN(n430) );
  INV_X4 U1032 ( .A(inputSRAM_Data[6]), .ZN(n431) );
  INV_X4 U1033 ( .A(inputSRAM_Data[5]), .ZN(n432) );
  INV_X4 U1034 ( .A(inputSRAM_Data[4]), .ZN(n433) );
  INV_X4 U1035 ( .A(inputSRAM_Data[3]), .ZN(n434) );
  INV_X4 U1039 ( .A(graphRead1_DataInput[71]), .ZN(n438) );
  INV_X4 U1040 ( .A(graphRead1_DataInput[70]), .ZN(n439) );
  INV_X4 U1041 ( .A(graphRead1_DataInput[69]), .ZN(n440) );
  INV_X4 U1042 ( .A(graphRead1_DataInput[68]), .ZN(n441) );
  INV_X4 U1043 ( .A(graphRead1_DataInput[67]), .ZN(n442) );
  INV_X4 U1044 ( .A(graphRead1_DataInput[66]), .ZN(n443) );
  INV_X4 U1045 ( .A(graphRead1_DataInput[65]), .ZN(n444) );
  INV_X4 U1046 ( .A(graphRead1_DataInput[64]), .ZN(n445) );
  INV_X4 U1049 ( .A(graphRead1_DataInput[10]), .ZN(n448) );
  INV_X4 U1050 ( .A(graphRead1_DataInput[9]), .ZN(n449) );
  INV_X4 U1051 ( .A(graphRead1_DataInput[8]), .ZN(n450) );
  INV_X4 U1052 ( .A(graphRead1_DataInput[7]), .ZN(n451) );
  INV_X4 U1053 ( .A(graphRead1_DataInput[6]), .ZN(n452) );
  INV_X4 U1054 ( .A(graphRead1_DataInput[5]), .ZN(n453) );
  INV_X4 U1055 ( .A(graphRead1_DataInput[4]), .ZN(n454) );
  INV_X4 U1056 ( .A(graphRead1_DataInput[3]), .ZN(n455) );
  INV_X4 U1057 ( .A(graphRead1_DataInput[2]), .ZN(n456) );
  INV_X4 U1060 ( .A(graphRead2_DataInput[127]), .ZN(n459) );
  INV_X4 U1061 ( .A(graphRead2_DataInput[126]), .ZN(n460) );
  INV_X4 U1062 ( .A(graphRead2_DataInput[125]), .ZN(n461) );
  INV_X4 U1063 ( .A(graphRead2_DataInput[124]), .ZN(n462) );
  INV_X4 U1064 ( .A(graphRead2_DataInput[123]), .ZN(n463) );
  INV_X4 U1065 ( .A(graphRead2_DataInput[122]), .ZN(n464) );
  INV_X4 U1066 ( .A(graphRead2_DataInput[121]), .ZN(n465) );
  INV_X4 U1067 ( .A(graphRead2_DataInput[120]), .ZN(n466) );
  INV_X4 U1068 ( .A(graphRead2_DataInput[119]), .ZN(n467) );
  INV_X4 U1069 ( .A(graphRead2_DataInput[118]), .ZN(n468) );
  INV_X4 U1070 ( .A(graphRead2_DataInput[117]), .ZN(n469) );
  INV_X4 U1071 ( .A(graphRead2_DataInput[116]), .ZN(n470) );
  INV_X4 U1072 ( .A(graphRead2_DataInput[115]), .ZN(n471) );
  INV_X4 U1073 ( .A(graphRead2_DataInput[114]), .ZN(n472) );
  INV_X4 U1074 ( .A(graphRead2_DataInput[113]), .ZN(n473) );
  INV_X4 U1075 ( .A(graphRead2_DataInput[112]), .ZN(n474) );
  INV_X4 U1076 ( .A(graphRead2_DataInput[111]), .ZN(n475) );
  INV_X4 U1077 ( .A(graphRead2_DataInput[110]), .ZN(n476) );
  INV_X4 U1078 ( .A(graphRead2_DataInput[109]), .ZN(n477) );
  INV_X4 U1079 ( .A(graphRead2_DataInput[108]), .ZN(n478) );
  INV_X4 U1080 ( .A(graphRead2_DataInput[107]), .ZN(n479) );
  INV_X4 U1081 ( .A(graphRead2_DataInput[106]), .ZN(n480) );
  INV_X4 U1082 ( .A(graphRead2_DataInput[105]), .ZN(n481) );
  INV_X4 U1083 ( .A(graphRead2_DataInput[104]), .ZN(n482) );
  INV_X4 U1084 ( .A(graphRead2_DataInput[95]), .ZN(n483) );
  INV_X4 U1085 ( .A(graphRead2_DataInput[94]), .ZN(n484) );
  INV_X4 U1086 ( .A(graphRead2_DataInput[93]), .ZN(n485) );
  INV_X4 U1087 ( .A(graphRead2_DataInput[92]), .ZN(n486) );
  INV_X4 U1088 ( .A(graphRead2_DataInput[91]), .ZN(n487) );
  INV_X4 U1089 ( .A(graphRead2_DataInput[90]), .ZN(n488) );
  INV_X4 U1090 ( .A(graphRead2_DataInput[89]), .ZN(n489) );
  INV_X4 U1091 ( .A(graphRead2_DataInput[88]), .ZN(n490) );
  INV_X4 U1092 ( .A(graphRead2_DataInput[87]), .ZN(n491) );
  INV_X4 U1093 ( .A(graphRead2_DataInput[86]), .ZN(n492) );
  INV_X4 U1100 ( .A(graphRead2_DataInput[79]), .ZN(n499) );
  INV_X4 U1101 ( .A(graphRead2_DataInput[78]), .ZN(n500) );
  INV_X4 U1102 ( .A(graphRead2_DataInput[77]), .ZN(n501) );
  INV_X4 U1103 ( .A(graphRead2_DataInput[76]), .ZN(n502) );
  INV_X4 U1104 ( .A(graphRead2_DataInput[75]), .ZN(n503) );
  INV_X4 U1105 ( .A(graphRead2_DataInput[74]), .ZN(n504) );
  INV_X4 U1106 ( .A(graphRead2_DataInput[73]), .ZN(n505) );
  INV_X4 U1107 ( .A(graphRead2_DataInput[72]), .ZN(n506) );
  INV_X4 U1108 ( .A(graphRead2_DataInput[71]), .ZN(n507) );
  INV_X4 U1109 ( .A(graphRead2_DataInput[70]), .ZN(n508) );
  INV_X4 U1116 ( .A(graphRead2_DataInput[63]), .ZN(n515) );
  INV_X4 U1117 ( .A(graphRead2_DataInput[62]), .ZN(n516) );
  INV_X4 U1118 ( .A(graphRead2_DataInput[61]), .ZN(n517) );
  INV_X4 U1119 ( .A(graphRead2_DataInput[60]), .ZN(n518) );
  INV_X4 U1120 ( .A(graphRead2_DataInput[59]), .ZN(n519) );
  INV_X4 U1121 ( .A(graphRead2_DataInput[58]), .ZN(n520) );
  INV_X4 U1122 ( .A(graphRead2_DataInput[57]), .ZN(n521) );
  INV_X4 U1123 ( .A(graphRead2_DataInput[56]), .ZN(n522) );
  INV_X4 U1124 ( .A(graphRead2_DataInput[47]), .ZN(n523) );
  INV_X4 U1125 ( .A(graphRead2_DataInput[46]), .ZN(n524) );
  INV_X4 U1126 ( .A(graphRead2_DataInput[45]), .ZN(n525) );
  INV_X4 U1127 ( .A(graphRead2_DataInput[44]), .ZN(n526) );
  INV_X4 U1128 ( .A(graphRead2_DataInput[43]), .ZN(n527) );
  INV_X4 U1129 ( .A(graphRead2_DataInput[42]), .ZN(n528) );
  INV_X4 U1130 ( .A(graphRead2_DataInput[41]), .ZN(n529) );
  INV_X4 U1131 ( .A(graphRead2_DataInput[40]), .ZN(n530) );
  INV_X4 U1132 ( .A(graphRead2_DataInput[31]), .ZN(n531) );
  INV_X4 U1133 ( .A(graphRead2_DataInput[30]), .ZN(n532) );
  INV_X4 U1134 ( .A(graphRead2_DataInput[29]), .ZN(n533) );
  INV_X4 U1135 ( .A(graphRead2_DataInput[28]), .ZN(n534) );
  INV_X4 U1136 ( .A(graphRead2_DataInput[27]), .ZN(n535) );
  INV_X4 U1137 ( .A(graphRead2_DataInput[26]), .ZN(n536) );
  INV_X4 U1138 ( .A(graphRead2_DataInput[25]), .ZN(n537) );
  INV_X4 U1139 ( .A(graphRead2_DataInput[24]), .ZN(n538) );
  INV_X4 U1140 ( .A(graphRead2_DataInput[23]), .ZN(n539) );
  INV_X4 U1141 ( .A(graphRead2_DataInput[22]), .ZN(n540) );
  INV_X4 U1148 ( .A(graphRead2_DataInput[15]), .ZN(n547) );
  INV_X4 U1149 ( .A(graphRead2_DataInput[14]), .ZN(n548) );
  INV_X4 U1150 ( .A(graphRead2_DataInput[13]), .ZN(n549) );
  INV_X4 U1151 ( .A(graphRead2_DataInput[12]), .ZN(n550) );
  INV_X4 U1152 ( .A(graphRead2_DataInput[11]), .ZN(n551) );
  INV_X4 U1153 ( .A(graphRead2_DataInput[10]), .ZN(n552) );
  INV_X4 U1154 ( .A(graphRead2_DataInput[9]), .ZN(n553) );
  INV_X4 U1155 ( .A(graphRead2_DataInput[8]), .ZN(n554) );
  INV_X4 U1156 ( .A(graphRead2_DataInput[7]), .ZN(n555) );
  INV_X4 U1157 ( .A(graphRead2_DataInput[6]), .ZN(n556) );
  INV_X4 U1164 ( .A(n1040), .ZN(n563) );
  INV_X4 U1165 ( .A(n845), .ZN(n564) );
  INV_X4 U1176 ( .A(state[1]), .ZN(n575) );
  OR2_X1 U1178 ( .A1(n637), .A2(n3157), .ZN(n577) );
  OR4_X1 U1193 ( .A1(n933), .A2(n934), .A3(n935), .A4(n936), .ZN(n932) );
  OR4_X1 U1194 ( .A1(n953), .A2(n954), .A3(n955), .A4(n956), .ZN(n931) );
  OR2_X1 U1195 ( .A1(graphRead1_DataInput[96]), .A2(graphRead1_DataInput[95]), 
        .ZN(n965) );
  AND2_X1 U1200 ( .A1(n1071), .A2(n1072), .ZN(graphData1_Zero_reg) );
  DFF_X2 offsetMux_Sel1_reg_1_ ( .D(n1377), .CK(clock), .Q(r572_A_1_), .QN(n60) );
  DFF_X2 offsetMux_Sel2_reg_0_ ( .D(n1287), .CK(clock), .Q(
        mult_add_378_aco_a_0_), .QN(n418) );
  DFF_X2 offsetMux_Sel2_reg_2_ ( .D(n1285), .CK(clock), .Q(
        mult_add_378_aco_a_2_), .QN(n416) );
  DFF_X2 offsetMux_Sel2_reg_1_ ( .D(n1286), .CK(clock), .Q(
        mult_add_378_aco_a_1_), .QN(n417) );
  DFF_X2 workWrite_Dist_reg_15_ ( .D(n1130), .CK(clock), .Q(workWrite_Dist[15]), .QN(n2921) );
  DFF_X2 iterStop_reg ( .D(n1154), .CK(clock), .Q(iterStop), .QN(n2813) );
  DFF_X2 workWrite_Dist_reg_14_ ( .D(n1131), .CK(clock), .Q(workWrite_Dist[14]), .QN(n2916) );
  DFF_X2 workWrite_Dist_reg_13_ ( .D(n1132), .CK(clock), .Q(workWrite_Dist[13]), .QN(n2913) );
  DFF_X2 workWrite_Dist_reg_11_ ( .D(n1134), .CK(clock), .Q(workWrite_Dist[11]) );
  DFF_X2 workWrite_Dist_reg_10_ ( .D(n1135), .CK(clock), .Q(workWrite_Dist[10]), .QN(n2905) );
  DFF_X2 workWrite_Dist_reg_8_ ( .D(n1137), .CK(clock), .Q(workWrite_Dist[8]), 
        .QN(n2896) );
  DFF_X2 workWrite_Dist_reg_6_ ( .D(n1139), .CK(clock), .Q(workWrite_Dist[6]), 
        .QN(net11164) );
  DFF_X2 workWrite_Dist_reg_1_ ( .D(n1144), .CK(clock), .Q(workWrite_Dist[1]), 
        .QN(n2873) );
  DFF_X2 workWrite_Dist_reg_12_ ( .D(n1133), .CK(clock), .Q(workWrite_Dist[12]), .QN(n2910) );
  DFF_X2 workWrite_Dist_reg_9_ ( .D(n1136), .CK(clock), .Q(workWrite_Dist[9]), 
        .QN(n2901) );
  DFF_X2 workWrite_Dist_reg_4_ ( .D(n1141), .CK(clock), .Q(workWrite_Dist[4]), 
        .QN(n2885) );
  DFF_X2 workWrite_Dist_reg_0_ ( .D(n1145), .CK(clock), .Q(workWrite_Dist[0]), 
        .QN(n2869) );
  DFF_X2 vertexCount_reg_3_ ( .D(n1331), .CK(clock), .Q(sub_387_A_3_), .QN(n39) );
  DFF_X2 vertexCount_reg_4_ ( .D(n1330), .CK(clock), .Q(sub_387_A_4_), .QN(n38) );
  DFF_X2 graphRead1_Addr_reg_1_ ( .D(n1349), .CK(clock), .Q(graphRead1_Addr[1]), .QN(n291) );
  DFF_X2 graphRead1_Addr_reg_2_ ( .D(n1348), .CK(clock), .Q(graphRead1_Addr[2]), .QN(n289) );
  DFF_X2 graphRead1_Addr_reg_3_ ( .D(n1347), .CK(clock), .Q(graphRead1_Addr[3]), .QN(n287) );
  DFF_X2 graphRead1_Addr_reg_4_ ( .D(n1346), .CK(clock), .Q(graphRead1_Addr[4]), .QN(n285) );
  DFF_X2 graphRead1_Addr_reg_5_ ( .D(n1345), .CK(clock), .Q(graphRead1_Addr[5]), .QN(n283) );
  DFF_X2 graphRead1_Addr_reg_6_ ( .D(n1344), .CK(clock), .Q(graphRead1_Addr[6]), .QN(n281) );
  DFF_X2 graphRead1_Addr_reg_7_ ( .D(n1343), .CK(clock), .Q(graphRead1_Addr[7]), .QN(n279) );
  DFF_X2 graphRead1_Addr_reg_0_ ( .D(n1350), .CK(clock), .Q(graphRead1_Addr[0]), .QN(n293) );
  DFF_X2 outputWrite_Addr_reg_0_ ( .D(n1321), .CK(clock), .Q(
        outputWrite_Addr[0]), .QN(n365) );
  XNOR2_X2 U119 ( .A(eq_565_B_1_), .B(U97_DATA2_1), .ZN(n668) );
  XNOR2_X2 U118 ( .A(eq_565_B_0_), .B(U97_DATA2_0), .ZN(n669) );
  XNOR2_X2 U121 ( .A(eq_565_B_3_), .B(U97_DATA2_3), .ZN(n666) );
  XNOR2_X2 U120 ( .A(eq_565_B_2_), .B(U97_DATA2_2), .ZN(n667) );
  XNOR2_X2 U114 ( .A(eq_565_B_5_), .B(U97_DATA2_5), .ZN(n664) );
  XNOR2_X2 U113 ( .A(eq_565_B_4_), .B(U97_DATA2_4), .ZN(n665) );
  XNOR2_X2 U116 ( .A(eq_565_B_7_), .B(U97_DATA2_7), .ZN(n662) );
  XNOR2_X2 U115 ( .A(eq_565_B_6_), .B(U97_DATA2_6), .ZN(n663) );
  DFF_X2 zeroFlag_reg ( .D(n71), .CK(clock), .Q(zeroFlag) );
  DFF_X2 workRead2_Dist_reg_14_ ( .D(n299), .CK(clock), .Q(U112_DATA1_14), 
        .QN(n2499) );
  DFF_X2 workRead2_Dist_reg_12_ ( .D(n301), .CK(clock), .Q(U112_DATA1_12), 
        .QN(n2488) );
  DFF_X2 workRead2_Dist_reg_10_ ( .D(n303), .CK(clock), .Q(U112_DATA1_10), 
        .QN(n2909) );
  DFF_X2 workRead2_Dist_reg_9_ ( .D(n304), .CK(clock), .Q(U112_DATA1_9), .QN(
        n2904) );
  DFF_X2 workRead2_Dist_reg_8_ ( .D(n305), .CK(clock), .Q(U112_DATA1_8), .QN(
        n2900) );
  DFF_X2 workRead2_Dist_reg_6_ ( .D(n307), .CK(clock), .Q(U112_DATA1_6), .QN(
        n2616) );
  DFF_X2 workRead2_Dist_reg_5_ ( .D(n308), .CK(clock), .Q(U112_DATA1_5), .QN(
        net11165) );
  DFF_X2 workRead2_Dist_reg_4_ ( .D(n309), .CK(clock), .Q(U112_DATA1_4), .QN(
        net11170) );
  DFF_X2 workRead2_Dist_reg_2_ ( .D(n311), .CK(clock), .Q(U112_DATA1_2), .QN(
        n2881) );
  DFF_X2 workRead2_Dist_reg_0_ ( .D(n313), .CK(clock), .Q(U112_DATA1_0), .QN(
        n2872) );
  DFF_X2 workRead2_Dist_reg_3_ ( .D(n310), .CK(clock), .Q(U112_DATA1_3), .QN(
        net11175) );
  DFF_X2 workRead1_Dist_reg_9_ ( .D(n1313), .CK(clock), .Q(U91_DATA2_1), .QN(
        n2474) );
  DFF_X2 workRead1_Dist_reg_8_ ( .D(n1312), .CK(clock), .Q(U91_DATA2_0), .QN(
        n2498) );
  DFF_X2 workRead1_Dist_reg_5_ ( .D(n1309), .CK(clock), .Q(U92_DATA2_5), .QN(
        n2481) );
  DFF_X2 graphRead2_Data_reg_112_ ( .D(n137), .CK(clock), .Q(U37_DATA1_0), 
        .QN(n2696) );
  DFF_X2 graphRead2_Data_reg_96_ ( .D(n154), .CK(clock), .Q(U37_DATA2_0), .QN(
        n2697) );
  DFF_X2 graphRead2_Data_reg_51_ ( .D(n199), .CK(clock), .Q(U37_DATA5_3), .QN(
        n2729) );
  DFF_X2 graphRead2_Data_reg_35_ ( .D(n215), .CK(clock), .Q(U37_DATA6_3), .QN(
        n2731) );
  DFF_X2 graphRead2_Data_reg_115_ ( .D(n131), .CK(clock), .Q(U37_DATA1_3), 
        .QN(n2724) );
  DFF_X2 graphRead2_Data_reg_114_ ( .D(n133), .CK(clock), .Q(U37_DATA1_2), 
        .QN(n2713) );
  DFF_X2 graphRead2_Data_reg_113_ ( .D(n135), .CK(clock), .Q(U37_DATA1_1), 
        .QN(net11592) );
  DFF_X2 graphRead2_Data_reg_99_ ( .D(n151), .CK(clock), .Q(U37_DATA2_3), .QN(
        n2725) );
  DFF_X2 graphRead2_Data_reg_98_ ( .D(n152), .CK(clock), .Q(U37_DATA2_2), .QN(
        n2714) );
  DFF_X2 graphRead2_Data_reg_97_ ( .D(n153), .CK(clock), .Q(U37_DATA2_1), .QN(
        net11590) );
  DFF_X2 graphRead2_Data_reg_50_ ( .D(n200), .CK(clock), .Q(U37_DATA5_2), .QN(
        n2718) );
  DFF_X2 graphRead2_Data_reg_49_ ( .D(n201), .CK(clock), .Q(U37_DATA5_1), .QN(
        net11586) );
  DFF_X2 graphRead2_Data_reg_48_ ( .D(n202), .CK(clock), .Q(U37_DATA5_0), .QN(
        n2701) );
  DFF_X2 graphRead2_Data_reg_34_ ( .D(n216), .CK(clock), .Q(U37_DATA6_2), .QN(
        n2720) );
  DFF_X2 graphRead2_Data_reg_33_ ( .D(n217), .CK(clock), .Q(U37_DATA6_1), .QN(
        net11584) );
  DFF_X2 graphRead2_Data_reg_32_ ( .D(n218), .CK(clock), .Q(U37_DATA6_0), .QN(
        n2703) );
  DFF_X2 graphRead2_Data_reg_119_ ( .D(n112), .CK(clock), .Q(U37_DATA1_7), 
        .QN(n2764) );
  DFF_X2 graphRead2_Data_reg_118_ ( .D(n125), .CK(clock), .Q(U37_DATA1_6), 
        .QN(n2757) );
  DFF_X2 graphRead2_Data_reg_117_ ( .D(n127), .CK(clock), .Q(U37_DATA1_5), 
        .QN(n2746) );
  DFF_X2 graphRead2_Data_reg_116_ ( .D(n129), .CK(clock), .Q(U37_DATA1_4), 
        .QN(n2735) );
  DFF_X2 graphRead2_Data_reg_102_ ( .D(n148), .CK(clock), .Q(U37_DATA2_6), 
        .QN(n2758) );
  DFF_X2 graphRead2_Data_reg_101_ ( .D(n149), .CK(clock), .Q(U37_DATA2_5), 
        .QN(n2747) );
  DFF_X2 graphRead2_Data_reg_100_ ( .D(n150), .CK(clock), .Q(U37_DATA2_4), 
        .QN(n2736) );
  DFF_X2 graphRead2_Data_reg_55_ ( .D(n195), .CK(clock), .Q(U37_DATA5_7), .QN(
        net11520) );
  DFF_X2 graphRead2_Data_reg_54_ ( .D(n196), .CK(clock), .Q(U37_DATA5_6), .QN(
        n2760) );
  DFF_X2 graphRead2_Data_reg_53_ ( .D(n197), .CK(clock), .Q(U37_DATA5_5), .QN(
        n2751) );
  DFF_X2 graphRead2_Data_reg_52_ ( .D(n198), .CK(clock), .Q(U37_DATA5_4), .QN(
        n2740) );
  DFF_X2 graphRead2_Data_reg_38_ ( .D(n212), .CK(clock), .Q(U37_DATA6_6), .QN(
        n2762) );
  DFF_X2 graphRead2_Data_reg_37_ ( .D(n213), .CK(clock), .Q(U37_DATA6_5), .QN(
        n2753) );
  DFF_X2 graphRead2_Data_reg_36_ ( .D(n214), .CK(clock), .Q(U37_DATA6_4), .QN(
        n2742) );
  DFF_X2 vertex_reg_7_ ( .D(n1374), .CK(clock), .Q(n2867), .QN(n62) );
  DFF_X2 vertex_reg_6_ ( .D(n1372), .CK(clock), .Q(n2864), .QN(n63) );
  DFF_X2 vertex_reg_5_ ( .D(n1370), .CK(clock), .Q(n2862), .QN(n64) );
  DFF_X2 vertex_reg_4_ ( .D(n1368), .CK(clock), .Q(n2860), .QN(n65) );
  DFF_X2 vertex_reg_3_ ( .D(n1366), .CK(clock), .Q(n2858), .QN(n66) );
  DFF_X2 vertex_reg_2_ ( .D(n1364), .CK(clock), .Q(n2856), .QN(n67) );
  DFF_X2 vertex_reg_1_ ( .D(n1362), .CK(clock), .Q(n2854), .QN(n68) );
  DFF_X2 vertex_reg_0_ ( .D(n1352), .CK(clock), .Q(n2852), .QN(n69) );
  DFF_X2 graphRead2_Data_reg_80_ ( .D(n1248), .CK(clock), .QN(n170) );
  DFF_X2 graphRead2_Data_reg_64_ ( .D(n1232), .CK(clock), .QN(n186) );
  DFF_X2 graphRead2_Data_reg_83_ ( .D(n1251), .CK(clock), .QN(n167) );
  DFF_X2 graphRead2_Data_reg_82_ ( .D(n1250), .CK(clock), .QN(n168) );
  DFF_X2 graphRead2_Data_reg_81_ ( .D(n1249), .CK(clock), .QN(n169) );
  DFF_X2 graphRead2_Data_reg_67_ ( .D(n1235), .CK(clock), .QN(n183) );
  DFF_X2 graphRead2_Data_reg_66_ ( .D(n1234), .CK(clock), .QN(n184) );
  DFF_X2 graphRead2_Data_reg_65_ ( .D(n1233), .CK(clock), .QN(n185) );
  DFF_X2 graphRead2_Data_reg_18_ ( .D(n1202), .CK(clock), .QN(n232) );
  DFF_X2 graphRead2_Data_reg_17_ ( .D(n1201), .CK(clock), .QN(n233) );
  DFF_X2 graphRead2_Data_reg_16_ ( .D(n1200), .CK(clock), .QN(n234) );
  DFF_X2 graphRead2_Data_reg_2_ ( .D(n1186), .CK(clock), .QN(n248) );
  DFF_X2 graphRead2_Data_reg_1_ ( .D(n1185), .CK(clock), .QN(n249) );
  DFF_X2 graphRead2_Data_reg_0_ ( .D(n1184), .CK(clock), .QN(n250) );
  DFF_X2 graphRead2_Data_reg_85_ ( .D(n1253), .CK(clock), .QN(n165) );
  DFF_X2 graphRead2_Data_reg_84_ ( .D(n1252), .CK(clock), .QN(n166) );
  DFF_X2 graphRead2_Data_reg_69_ ( .D(n1237), .CK(clock), .QN(n181) );
  DFF_X2 graphRead2_Data_reg_68_ ( .D(n1236), .CK(clock), .QN(n182) );
  DFF_X2 graphRead2_Data_reg_21_ ( .D(n1205), .CK(clock), .QN(n229) );
  DFF_X2 graphRead2_Data_reg_20_ ( .D(n1204), .CK(clock), .QN(n230) );
  DFF_X2 graphRead2_Data_reg_19_ ( .D(n1203), .CK(clock), .QN(n231) );
  DFF_X2 graphRead2_Data_reg_5_ ( .D(n1189), .CK(clock), .QN(n245) );
  DFF_X2 graphRead2_Data_reg_4_ ( .D(n1188), .CK(clock), .QN(n246) );
  DFF_X2 graphRead2_Data_reg_3_ ( .D(n1187), .CK(clock), .QN(n247) );
  DFF_X2 daughterCount_reg_4_ ( .D(n1400), .CK(clock), .QN(n333) );
  DFF_X2 daughterCount_reg_3_ ( .D(n1401), .CK(clock), .QN(n334) );
  DFF_X2 daughterCount_reg_2_ ( .D(n1402), .CK(clock), .QN(n335) );
  DFF_X2 graphRead2_Data_reg_31_ ( .D(n1215), .CK(clock), .QN(n219) );
  DFF_X2 graphRead2_Data_reg_30_ ( .D(n1214), .CK(clock), .QN(n220) );
  DFF_X2 graphRead2_Data_reg_29_ ( .D(n1213), .CK(clock), .QN(n221) );
  DFF_X2 graphRead2_Data_reg_15_ ( .D(n1199), .CK(clock), .QN(n235) );
  DFF_X2 graphRead2_Data_reg_14_ ( .D(n1198), .CK(clock), .QN(n236) );
  DFF_X2 graphRead2_Data_reg_13_ ( .D(n1197), .CK(clock), .QN(n237) );
  DFF_X2 graphRead2_Data_reg_28_ ( .D(n1212), .CK(clock), .QN(n222) );
  DFF_X2 graphRead2_Data_reg_27_ ( .D(n1211), .CK(clock), .QN(n223) );
  DFF_X2 graphRead2_Data_reg_26_ ( .D(n1210), .CK(clock), .QN(n224) );
  DFF_X2 graphRead2_Data_reg_25_ ( .D(n1209), .CK(clock), .QN(n225) );
  DFF_X2 graphRead2_Data_reg_24_ ( .D(n1208), .CK(clock), .QN(n226) );
  DFF_X2 graphRead2_Data_reg_12_ ( .D(n1196), .CK(clock), .QN(n238) );
  DFF_X2 graphRead2_Data_reg_11_ ( .D(n1195), .CK(clock), .QN(n239) );
  DFF_X2 graphRead2_Data_reg_10_ ( .D(n1194), .CK(clock), .QN(n240) );
  DFF_X2 graphRead2_Data_reg_9_ ( .D(n1193), .CK(clock), .QN(n241) );
  DFF_X2 graphRead2_Data_reg_8_ ( .D(n1192), .CK(clock), .QN(n242) );
  DFF_X2 graphRead2_Data_reg_87_ ( .D(n1255), .CK(clock), .QN(n163) );
  DFF_X2 graphRead2_Data_reg_71_ ( .D(n1239), .CK(clock), .QN(n179) );
  DFF_X2 graphRead2_Data_reg_22_ ( .D(n1206), .CK(clock), .QN(n228) );
  DFF_X2 graphRead2_Data_reg_7_ ( .D(n1191), .CK(clock), .Q(n2596), .QN(n243)
         );
  DFF_X2 graphRead2_Data_reg_6_ ( .D(n1190), .CK(clock), .QN(n244) );
  DFF_X2 graphRead2_Data_reg_86_ ( .D(n1254), .CK(clock), .QN(n164) );
  DFF_X2 graphRead2_Data_reg_70_ ( .D(n1238), .CK(clock), .QN(n180) );
  DFF_X2 graphRead2_Data_reg_23_ ( .D(n1207), .CK(clock), .QN(n227) );
  DFF_X2 totalVertex_reg_7_ ( .D(n1335), .CK(clock), .QN(n80) );
  DFF_X2 totalVertex_reg_6_ ( .D(n1336), .CK(clock), .QN(n81) );
  DFF_X2 totalVertex_reg_5_ ( .D(n1337), .CK(clock), .QN(n82) );
  DFF_X2 totalVertex_reg_4_ ( .D(n1338), .CK(clock), .QN(n83) );
  DFF_X2 totalVertex_reg_3_ ( .D(n1339), .CK(clock), .QN(n84) );
  DFF_X2 totalVertex_reg_2_ ( .D(n1340), .CK(clock), .QN(n85) );
  DFF_X2 workRead1_Pred_reg_7_ ( .D(n1386), .CK(clock), .Q(U97_DATA4_7), .QN(
        n2) );
  DFF_X2 workRead1_Pred_reg_6_ ( .D(n1385), .CK(clock), .Q(U97_DATA4_6), .QN(
        n3) );
  DFF_X2 workRead1_Pred_reg_5_ ( .D(n1384), .CK(clock), .Q(U97_DATA4_5), .QN(
        n4) );
  DFF_X2 workRead1_Pred_reg_4_ ( .D(n1383), .CK(clock), .Q(U97_DATA4_4), .QN(
        n5) );
  DFF_X2 workRead1_Pred_reg_3_ ( .D(n1382), .CK(clock), .Q(U97_DATA4_3), .QN(
        n6) );
  DFF_X2 workRead1_Pred_reg_2_ ( .D(n1381), .CK(clock), .Q(U97_DATA4_2), .QN(
        n7) );
  DFF_X2 workRead1_Pred_reg_1_ ( .D(n1380), .CK(clock), .Q(U97_DATA4_1), .QN(
        n8) );
  DFF_X2 workRead1_Pred_reg_0_ ( .D(n1379), .CK(clock), .Q(U97_DATA4_0), .QN(
        n9) );
  DFF_X2 destReg_reg_3_ ( .D(n1417), .CK(clock), .Q(U97_DATA3_3), .QN(n3104)
         );
  DFF_X2 destReg_reg_5_ ( .D(n1419), .CK(clock), .Q(U97_DATA3_5), .QN(n3108)
         );
  DFF_X2 destReg_reg_4_ ( .D(n1418), .CK(clock), .Q(U97_DATA3_4), .QN(n3106)
         );
  DFF_X2 destReg_reg_6_ ( .D(n1420), .CK(clock), .Q(U97_DATA3_6), .QN(n3110)
         );
  DFF_X2 destReg_reg_7_ ( .D(n1421), .CK(clock), .Q(U97_DATA3_7), .QN(n3112)
         );
  DFF_X2 destReg_reg_2_ ( .D(n1416), .CK(clock), .QN(n3102) );
  DFF_X2 destReg_reg_1_ ( .D(n1415), .CK(clock), .QN(n3100) );
  DFF_X2 destReg_reg_0_ ( .D(n1414), .CK(clock), .QN(n3098) );
  DFF_X2 sourceReg_reg_5_ ( .D(n1410), .CK(clock), .Q(eq_565_B_5_), .QN(n90)
         );
  DFF_X2 sourceReg_reg_4_ ( .D(n1409), .CK(clock), .Q(eq_565_B_4_), .QN(n91)
         );
  DFF_X2 sourceReg_reg_3_ ( .D(n1408), .CK(clock), .Q(eq_565_B_3_), .QN(n92)
         );
  DFF_X2 sourceReg_reg_7_ ( .D(n1412), .CK(clock), .Q(eq_565_B_7_), .QN(n88)
         );
  DFF_X2 sourceReg_reg_6_ ( .D(n1411), .CK(clock), .Q(eq_565_B_6_), .QN(n89)
         );
  DFF_X2 sourceReg_reg_2_ ( .D(n1407), .CK(clock), .Q(eq_565_B_2_), .QN(n93)
         );
  DFF_X2 sourceReg_reg_1_ ( .D(n1406), .CK(clock), .Q(eq_565_B_1_), .QN(n94)
         );
  DFF_X2 sourceReg_reg_0_ ( .D(n1405), .CK(clock), .Q(eq_565_B_0_), .QN(n95)
         );
  DFF_X2 workRead2_Dist_reg_16_ ( .D(n297), .CK(clock), .Q(U112_DATA1_16), 
        .QN(n2484) );
  DFF_X2 workRead2_Dist_reg_15_ ( .D(n298), .CK(clock), .Q(U112_DATA1_15), 
        .QN(n2485) );
  DFF_X2 workRead2_Dist_reg_13_ ( .D(n300), .CK(clock), .Q(U112_DATA1_13), 
        .QN(n2486) );
  DFF_X2 workRead2_Dist_reg_11_ ( .D(n302), .CK(clock), .Q(U112_DATA1_11), 
        .QN(n2489) );
  DFF_X2 workRead2_Dist_reg_7_ ( .D(n306), .CK(clock), .Q(U112_DATA1_7), .QN(
        n2895) );
  DFF_X2 workRead2_Pred_reg_7_ ( .D(n314), .CK(clock), .Q(U113_DATA2_7), .QN(
        n391) );
  DFF_X2 workRead2_Pred_reg_6_ ( .D(n315), .CK(clock), .Q(U113_DATA2_6), .QN(
        n392) );
  DFF_X2 workRead2_Pred_reg_5_ ( .D(n316), .CK(clock), .Q(U113_DATA2_5), .QN(
        n393) );
  DFF_X2 workRead2_Pred_reg_4_ ( .D(n317), .CK(clock), .Q(U113_DATA2_4), .QN(
        n394) );
  DFF_X2 workRead2_Pred_reg_3_ ( .D(n318), .CK(clock), .Q(U113_DATA2_3), .QN(
        n395) );
  DFF_X2 workRead2_Pred_reg_2_ ( .D(n319), .CK(clock), .Q(U113_DATA2_2), .QN(
        n396) );
  DFF_X2 workRead2_Pred_reg_1_ ( .D(n320), .CK(clock), .Q(U113_DATA2_1), .QN(
        n397) );
  DFF_X2 workRead2_Pred_reg_0_ ( .D(n321), .CK(clock), .Q(U113_DATA2_0), .QN(
        n398) );
  DFF_X2 workRead2_Dist_reg_1_ ( .D(n312), .CK(clock), .Q(U112_DATA1_1), .QN(
        n2876) );
  DFF_X2 daughterCount_reg_1_ ( .D(n1403), .CK(clock), .Q(U3_U6_DATA4_1), .QN(
        n336) );
  DFF_X2 daughterCount_reg_5_ ( .D(n1399), .CK(clock), .Q(U3_U6_DATA4_5), .QN(
        n332) );
  DFF_X2 daughterCount_reg_6_ ( .D(n1398), .CK(clock), .Q(U3_U6_DATA4_6), .QN(
        n331) );
  DFF_X2 graphRead2_Data_reg_127_ ( .D(n1183), .CK(clock), .Q(U38_DATA1_7), 
        .QN(n104) );
  DFF_X2 graphRead2_Data_reg_126_ ( .D(n1182), .CK(clock), .Q(U38_DATA1_6), 
        .QN(n105) );
  DFF_X2 graphRead2_Data_reg_125_ ( .D(n1181), .CK(clock), .Q(U38_DATA1_5), 
        .QN(n106) );
  DFF_X2 graphRead2_Data_reg_111_ ( .D(n1175), .CK(clock), .Q(U38_DATA2_7), 
        .QN(n139) );
  DFF_X2 graphRead2_Data_reg_110_ ( .D(n1174), .CK(clock), .Q(U38_DATA2_6), 
        .QN(n140) );
  DFF_X2 graphRead2_Data_reg_109_ ( .D(n1173), .CK(clock), .Q(U38_DATA2_5), 
        .QN(n141) );
  DFF_X2 graphRead2_Data_reg_63_ ( .D(n1231), .CK(clock), .Q(U38_DATA5_7), 
        .QN(n187) );
  DFF_X2 graphRead2_Data_reg_62_ ( .D(n1230), .CK(clock), .Q(U38_DATA5_6), 
        .QN(n188) );
  DFF_X2 graphRead2_Data_reg_61_ ( .D(n1229), .CK(clock), .Q(U38_DATA5_5), 
        .QN(n189) );
  DFF_X2 graphRead2_Data_reg_46_ ( .D(n1222), .CK(clock), .Q(U38_DATA6_6), 
        .QN(n204) );
  DFF_X2 graphRead2_Data_reg_45_ ( .D(n1221), .CK(clock), .Q(U38_DATA6_5), 
        .QN(n205) );
  DFF_X2 graphRead2_Data_reg_44_ ( .D(n1220), .CK(clock), .Q(U38_DATA6_4), 
        .QN(n206) );
  DFF_X2 graphRead2_Data_reg_95_ ( .D(n1167), .CK(clock), .Q(U38_DATA3_7), 
        .QN(n155) );
  DFF_X2 graphRead2_Data_reg_94_ ( .D(n1166), .CK(clock), .Q(U38_DATA3_6), 
        .QN(n156) );
  DFF_X2 graphRead2_Data_reg_93_ ( .D(n1165), .CK(clock), .Q(U38_DATA3_5), 
        .QN(n157) );
  DFF_X2 graphRead2_Data_reg_79_ ( .D(n1247), .CK(clock), .Q(U38_DATA4_7), 
        .QN(n171) );
  DFF_X2 graphRead2_Data_reg_78_ ( .D(n1246), .CK(clock), .Q(U38_DATA4_6), 
        .QN(n172) );
  DFF_X2 graphRead2_Data_reg_77_ ( .D(n1245), .CK(clock), .Q(U38_DATA4_5), 
        .QN(n173) );
  DFF_X2 graphRead2_Data_reg_104_ ( .D(n1168), .CK(clock), .Q(U38_DATA2_0), 
        .QN(n146) );
  DFF_X2 graphRead2_Data_reg_47_ ( .D(n1223), .CK(clock), .Q(U38_DATA6_7), 
        .QN(n203) );
  DFF_X2 graphRead2_Data_reg_88_ ( .D(n1256), .CK(clock), .Q(U38_DATA3_0), 
        .QN(n162) );
  DFF_X2 graphRead2_Data_reg_72_ ( .D(n1240), .CK(clock), .Q(U38_DATA4_0), 
        .QN(n178) );
  DFF_X2 graphRead2_Data_reg_124_ ( .D(n1180), .CK(clock), .Q(U38_DATA1_4), 
        .QN(n107) );
  DFF_X2 graphRead2_Data_reg_123_ ( .D(n1179), .CK(clock), .Q(U38_DATA1_3), 
        .QN(n108) );
  DFF_X2 graphRead2_Data_reg_122_ ( .D(n1178), .CK(clock), .Q(U38_DATA1_2), 
        .QN(n109) );
  DFF_X2 graphRead2_Data_reg_121_ ( .D(n1177), .CK(clock), .Q(U38_DATA1_1), 
        .QN(n110) );
  DFF_X2 graphRead2_Data_reg_120_ ( .D(n1176), .CK(clock), .Q(U38_DATA1_0), 
        .QN(n111) );
  DFF_X2 graphRead2_Data_reg_108_ ( .D(n1172), .CK(clock), .Q(U38_DATA2_4), 
        .QN(n142) );
  DFF_X2 graphRead2_Data_reg_107_ ( .D(n1171), .CK(clock), .Q(U38_DATA2_3), 
        .QN(n143) );
  DFF_X2 graphRead2_Data_reg_106_ ( .D(n1170), .CK(clock), .Q(U38_DATA2_2), 
        .QN(n144) );
  DFF_X2 graphRead2_Data_reg_105_ ( .D(n1169), .CK(clock), .Q(U38_DATA2_1), 
        .QN(n145) );
  DFF_X2 graphRead2_Data_reg_60_ ( .D(n1228), .CK(clock), .Q(U38_DATA5_4), 
        .QN(n190) );
  DFF_X2 graphRead2_Data_reg_59_ ( .D(n1227), .CK(clock), .Q(U38_DATA5_3), 
        .QN(n191) );
  DFF_X2 graphRead2_Data_reg_58_ ( .D(n1226), .CK(clock), .Q(U38_DATA5_2), 
        .QN(n192) );
  DFF_X2 graphRead2_Data_reg_57_ ( .D(n1225), .CK(clock), .Q(U38_DATA5_1), 
        .QN(n193) );
  DFF_X2 graphRead2_Data_reg_56_ ( .D(n1224), .CK(clock), .Q(U38_DATA5_0), 
        .QN(n194) );
  DFF_X2 graphRead2_Data_reg_43_ ( .D(n1219), .CK(clock), .Q(U38_DATA6_3), 
        .QN(n207) );
  DFF_X2 graphRead2_Data_reg_42_ ( .D(n1218), .CK(clock), .Q(U38_DATA6_2), 
        .QN(n208) );
  DFF_X2 graphRead2_Data_reg_41_ ( .D(n1217), .CK(clock), .Q(U38_DATA6_1), 
        .QN(n209) );
  DFF_X2 graphRead2_Data_reg_40_ ( .D(n1216), .CK(clock), .Q(U38_DATA6_0), 
        .QN(n210) );
  DFF_X2 graphRead2_Data_reg_92_ ( .D(n1164), .CK(clock), .Q(U38_DATA3_4), 
        .QN(n158) );
  DFF_X2 graphRead2_Data_reg_91_ ( .D(n1163), .CK(clock), .Q(U38_DATA3_3), 
        .QN(n159) );
  DFF_X2 graphRead2_Data_reg_90_ ( .D(n1258), .CK(clock), .Q(U38_DATA3_2), 
        .QN(n160) );
  DFF_X2 graphRead2_Data_reg_89_ ( .D(n1257), .CK(clock), .Q(U38_DATA3_1), 
        .QN(n161) );
  DFF_X2 graphRead2_Data_reg_76_ ( .D(n1244), .CK(clock), .Q(U38_DATA4_4), 
        .QN(n174) );
  DFF_X2 graphRead2_Data_reg_75_ ( .D(n1243), .CK(clock), .Q(U38_DATA4_3), 
        .QN(n175) );
  DFF_X2 graphRead2_Data_reg_74_ ( .D(n1242), .CK(clock), .Q(U38_DATA4_2), 
        .QN(n176) );
  DFF_X2 graphRead2_Data_reg_73_ ( .D(n1241), .CK(clock), .Q(U38_DATA4_1), 
        .QN(n177) );
  DFF_X2 offsetMux_Sel1_reg_0_ ( .D(n1378), .CK(clock), .Q(r572_A_0_), .QN(n61) );
  DFF_X2 offsetMux_Sel1_reg_2_ ( .D(n1376), .CK(clock), .Q(r572_A_2_), .QN(n59) );
  DFF_X2 vertexNumber_reg_7_ ( .D(n1375), .CK(clock), .Q(U97_DATA2_7), .QN(n43) );
  DFF_X2 vertexNumber_reg_6_ ( .D(n1373), .CK(clock), .Q(U97_DATA2_6), .QN(n47) );
  DFF_X2 vertexNumber_reg_5_ ( .D(n1371), .CK(clock), .Q(U97_DATA2_5), .QN(n48) );
  DFF_X2 vertexNumber_reg_4_ ( .D(n1369), .CK(clock), .Q(U97_DATA2_4), .QN(n49) );
  DFF_X2 vertexNumber_reg_3_ ( .D(n1367), .CK(clock), .Q(U97_DATA2_3), .QN(n50) );
  DFF_X2 vertexNumber_reg_2_ ( .D(n1365), .CK(clock), .Q(U97_DATA2_2), .QN(n51) );
  DFF_X2 vertexNumber_reg_1_ ( .D(n1363), .CK(clock), .Q(U97_DATA2_1), .QN(n52) );
  DFF_X2 vertexNumber_reg_0_ ( .D(n1361), .CK(clock), .Q(U97_DATA2_0), .QN(n53) );
  DFF_X2 daughterCount_reg_7_ ( .D(n1397), .CK(clock), .Q(U3_U6_DATA4_7), .QN(
        n294) );
  DFF_X2 workWrite_Dist_reg_7_ ( .D(n1138), .CK(clock), .Q(workWrite_Dist[7]), 
        .QN(n2891) );
  DFF_X2 workWrite_Dist_reg_5_ ( .D(n1140), .CK(clock), .Q(workWrite_Dist[5]), 
        .QN(n2888) );
  DFF_X2 workWrite_Dist_reg_3_ ( .D(n1142), .CK(clock), .Q(workWrite_Dist[3]), 
        .QN(n2882) );
  DFF_X2 workWrite_Dist_reg_2_ ( .D(n1143), .CK(clock), .Q(workWrite_Dist[2]), 
        .QN(n2877) );
  DFF_X2 workWrite_Addr_reg_5_ ( .D(n1123), .CK(clock), .Q(workWrite_Addr[5]), 
        .QN(n2463) );
  DFF_X2 workWrite_Addr_reg_4_ ( .D(n1124), .CK(clock), .Q(workWrite_Addr[4]), 
        .QN(n2445) );
  DFF_X2 workWrite_Addr_reg_3_ ( .D(n1125), .CK(clock), .Q(workWrite_Addr[3]), 
        .QN(n2440) );
  DFF_X2 workWrite_Addr_reg_2_ ( .D(n1126), .CK(clock), .Q(workWrite_Addr[2]), 
        .QN(n2438) );
  DFF_X2 workWrite_Addr_reg_1_ ( .D(n1127), .CK(clock), .Q(workWrite_Addr[1]), 
        .QN(n2435) );
  DFF_X2 workWrite_Addr_reg_0_ ( .D(n1128), .CK(clock), .Q(workWrite_Addr[0]), 
        .QN(n2432) );
  DFF_X2 workRead1_Dist_reg_11_ ( .D(n1315), .CK(clock), .Q(U91_DATA2_3), .QN(
        n2495) );
  DFF_X2 workRead1_Dist_reg_15_ ( .D(n1319), .CK(clock), .Q(U91_DATA2_7), .QN(
        n2494) );
  DFF_X2 workRead1_Dist_reg_6_ ( .D(n1310), .CK(clock), .Q(U92_DATA2_6), .QN(
        n2493) );
  DFF_X2 workRead1_Dist_reg_13_ ( .D(n1317), .CK(clock), .Q(U91_DATA2_5), .QN(
        n2497) );
  DFF_X2 workRead1_Dist_reg_12_ ( .D(n1316), .CK(clock), .Q(U91_DATA2_4), .QN(
        n2492) );
  DFF_X2 workRead1_Dist_reg_10_ ( .D(n1314), .CK(clock), .Q(U91_DATA2_2), .QN(
        n2491) );
  DFF_X2 workRead1_Dist_reg_4_ ( .D(n1308), .CK(clock), .Q(U92_DATA2_4), .QN(
        n2490) );
  DFF_X2 workWrite_Addr_reg_7_ ( .D(n1121), .CK(clock), .Q(workWrite_Addr[7])
         );
  DFF_X2 workWrite_Addr_reg_6_ ( .D(n1122), .CK(clock), .Q(workWrite_Addr[6])
         );
  DFF_X2 outputWrite_Addr_reg_13_ ( .D(n351), .CK(clock), .Q(
        outputWrite_Addr[13]), .QN(n2453) );
  DFF_X2 outputWrite_Addr_reg_12_ ( .D(n363), .CK(clock), .Q(
        outputWrite_Addr[12]), .QN(n2468) );
  DFF_X2 outputWrite_Addr_reg_11_ ( .D(n362), .CK(clock), .Q(
        outputWrite_Addr[11]), .QN(n2462) );
  DFF_X2 outputWrite_Addr_reg_10_ ( .D(n361), .CK(clock), .Q(
        outputWrite_Addr[10]), .QN(n2456) );
  DFF_X2 outputWrite_Addr_reg_9_ ( .D(n360), .CK(clock), .Q(
        outputWrite_Addr[9]), .QN(n2466) );
  DFF_X2 outputWrite_Addr_reg_8_ ( .D(n359), .CK(clock), .Q(
        outputWrite_Addr[8]), .QN(n2461) );
  DFF_X2 outputWrite_Addr_reg_7_ ( .D(n358), .CK(clock), .Q(
        outputWrite_Addr[7]), .QN(n2449) );
  DFF_X2 outputWrite_Addr_reg_6_ ( .D(n357), .CK(clock), .Q(
        outputWrite_Addr[6]), .QN(n2465) );
  DFF_X2 outputWrite_Addr_reg_5_ ( .D(n356), .CK(clock), .Q(
        outputWrite_Addr[5]), .QN(n2460) );
  DFF_X2 outputWrite_Addr_reg_4_ ( .D(n355), .CK(clock), .Q(
        outputWrite_Addr[4]), .QN(n2455) );
  DFF_X2 outputWrite_Addr_reg_3_ ( .D(n354), .CK(clock), .Q(
        outputWrite_Addr[3]), .QN(n2464) );
  DFF_X2 outputWrite_Addr_reg_2_ ( .D(n353), .CK(clock), .Q(
        outputWrite_Addr[2]), .QN(n2459) );
  DFF_X2 outputWrite_Addr_reg_1_ ( .D(n352), .CK(clock), .Q(
        outputWrite_Addr[1]), .QN(n2454) );
  DFF_X2 graphRead2_Data_reg_39_ ( .D(n211), .CK(clock), .Q(U37_DATA6_7), .QN(
        net11518) );
  DFF_X2 graphRead2_Data_reg_103_ ( .D(n147), .CK(clock), .Q(U37_DATA2_7), 
        .QN(n2765) );
  DFF_X2 workRead1_Addr_reg_7_ ( .D(n1353), .CK(clock), .Q(workRead1_Addr[7]), 
        .QN(n2457) );
  DFF_X2 workRead1_Addr_reg_6_ ( .D(n1354), .CK(clock), .Q(workRead1_Addr[6]), 
        .QN(n2450) );
  DFF_X2 workRead1_Addr_reg_5_ ( .D(n1355), .CK(clock), .Q(workRead1_Addr[5]), 
        .QN(n2447) );
  DFF_X2 workRead1_Addr_reg_4_ ( .D(n1356), .CK(clock), .Q(workRead1_Addr[4]), 
        .QN(n2439) );
  DFF_X2 workRead1_Addr_reg_3_ ( .D(n1357), .CK(clock), .Q(workRead1_Addr[3]), 
        .QN(n2444) );
  DFF_X2 workRead1_Addr_reg_2_ ( .D(n1358), .CK(clock), .Q(workRead1_Addr[2]), 
        .QN(n2434) );
  DFF_X2 workRead1_Addr_reg_1_ ( .D(n1359), .CK(clock), .Q(workRead1_Addr[1]), 
        .QN(n2437) );
  DFF_X2 workRead1_Addr_reg_0_ ( .D(n1360), .CK(clock), .Q(workRead1_Addr[0])
         );
  DFF_X2 output_WE_reg ( .D(n1413), .CK(clock), .Q(output_WE) );
  DFF_X2 work_WE_reg ( .D(n1351), .CK(clock), .Q(work_WE) );
  DFF_X2 workWrite_Pred_reg_5_ ( .D(n1148), .CK(clock), .Q(workWrite_Pred[5])
         );
  DFF_X2 workWrite_Pred_reg_3_ ( .D(n1150), .CK(clock), .Q(workWrite_Pred[3])
         );
  DFF_X2 workWrite_Pred_reg_2_ ( .D(n1151), .CK(clock), .Q(workWrite_Pred[2])
         );
  DFF_X2 workWrite_Pred_reg_0_ ( .D(n1153), .CK(clock), .Q(workWrite_Pred[0])
         );
  DFF_X2 workWrite_Dist_reg_16_ ( .D(n1129), .CK(clock), .Q(workWrite_Dist[16]) );
  DFF_X2 vertexCount_reg_0_ ( .D(n1334), .CK(clock), .Q(sub_387_A_0_), .QN(
        n2467) );
  DFF_X2 workWrite_Pred_reg_7_ ( .D(n1146), .CK(clock), .Q(workWrite_Pred[7])
         );
  DFF_X2 workWrite_Pred_reg_6_ ( .D(n1147), .CK(clock), .Q(workWrite_Pred[6])
         );
  DFF_X2 workWrite_Pred_reg_4_ ( .D(n1149), .CK(clock), .Q(workWrite_Pred[4])
         );
  DFF_X2 workWrite_Pred_reg_1_ ( .D(n1152), .CK(clock), .Q(workWrite_Pred[1])
         );
  OAI22_X2 U692 ( .A1(n1041), .A2(n252), .B1(n1042), .B2(n251), .ZN(n1387) );
  NOR2_X2 U868 ( .A1(state[3]), .A2(state[2]), .ZN(n1054) );
  INV_X4 U18 ( .A(1'b1), .ZN(workWrite_Addr[8]) );
  INV_X4 U21 ( .A(1'b1), .ZN(workWrite_Addr[9]) );
  INV_X4 U23 ( .A(1'b1), .ZN(workWrite_Addr[10]) );
  INV_X4 U25 ( .A(1'b1), .ZN(workWrite_Addr[11]) );
  INV_X4 U28 ( .A(1'b1), .ZN(workWrite_Addr[12]) );
  INV_X4 U30 ( .A(1'b1), .ZN(workRead2_Addr[8]) );
  INV_X4 U32 ( .A(1'b1), .ZN(workRead2_Addr[9]) );
  INV_X4 U34 ( .A(1'b1), .ZN(workRead2_Addr[10]) );
  INV_X4 U36 ( .A(1'b1), .ZN(workRead2_Addr[11]) );
  INV_X4 U38 ( .A(1'b1), .ZN(workRead2_Addr[12]) );
  INV_X4 U40 ( .A(1'b1), .ZN(workRead1_Addr[8]) );
  INV_X4 U42 ( .A(1'b1), .ZN(workRead1_Addr[9]) );
  INV_X4 U44 ( .A(1'b1), .ZN(workRead1_Addr[10]) );
  INV_X4 U46 ( .A(1'b1), .ZN(workRead1_Addr[11]) );
  INV_X4 U48 ( .A(1'b1), .ZN(workRead1_Addr[12]) );
  AND2_X2 U50 ( .A1(mult_add_378_aco_a_0_), .A2(n2626), .ZN(n2482) );
  NAND2_X2 U51 ( .A1(net12979), .A2(net10884), .ZN(n2470) );
  NAND2_X4 U52 ( .A1(net12979), .A2(net10884), .ZN(net11742) );
  OAI221_X1 U53 ( .B1(n2484), .B2(net11742), .C1(n2483), .C2(net11750), .A(
        n2922), .ZN(n1129) );
  OAI221_X1 U54 ( .B1(n392), .B2(net11742), .C1(n63), .C2(net11894), .A(n2865), 
        .ZN(n1147) );
  OAI221_X1 U55 ( .B1(n395), .B2(n2470), .C1(n66), .C2(net11750), .A(n2859), 
        .ZN(n1150) );
  OAI221_X1 U56 ( .B1(n398), .B2(net11742), .C1(n69), .C2(net11894), .A(n2853), 
        .ZN(n1153) );
  OAI221_X1 U57 ( .B1(n394), .B2(net11742), .C1(n65), .C2(net11750), .A(n2861), 
        .ZN(n1149) );
  OAI221_X1 U58 ( .B1(n397), .B2(n2470), .C1(n68), .C2(net11750), .A(n2855), 
        .ZN(n1152) );
  NAND2_X4 U59 ( .A1(n2561), .A2(net13049), .ZN(net10761) );
  AOI22_X2 U60 ( .A1(net11466), .A2(U92_DATA2_2), .B1(net13034), .B2(net12622), 
        .ZN(net12620) );
  OAI21_X2 U61 ( .B1(net15569), .B2(n2564), .A(n2575), .ZN(n2593) );
  AOI21_X2 U62 ( .B1(n2549), .B2(U112_DATA1_16), .A(n2479), .ZN(n2515) );
  OAI221_X2 U63 ( .B1(n2432), .B2(n3116), .C1(n577), .C2(n53), .A(n630), .ZN(
        n1128) );
  OAI222_X2 U64 ( .A1(n2433), .A2(n265), .B1(n335), .B2(n3068), .C1(n472), 
        .C2(n2565), .ZN(n1402) );
  INV_X4 U65 ( .A(n2573), .ZN(n2433) );
  OAI21_X2 U66 ( .B1(n2549), .B2(U112_DATA1_16), .A(n2550), .ZN(n2514) );
  OAI22_X2 U67 ( .A1(n2434), .A2(n54), .B1(n1001), .B2(n989), .ZN(n1358) );
  OAI221_X2 U68 ( .B1(n2435), .B2(n3116), .C1(n577), .C2(n52), .A(n624), .ZN(
        n1127) );
  OAI222_X2 U69 ( .A1(n2436), .A2(n263), .B1(n334), .B2(n3068), .C1(n471), 
        .C2(n2565), .ZN(n1401) );
  INV_X4 U70 ( .A(n2573), .ZN(n2436) );
  OAI22_X2 U71 ( .A1(n2437), .A2(n54), .B1(n1003), .B2(n989), .ZN(n1359) );
  OAI221_X2 U72 ( .B1(n2438), .B2(n3116), .C1(n577), .C2(n51), .A(n618), .ZN(
        n1126) );
  OAI221_X1 U73 ( .B1(n2872), .B2(n2470), .C1(n2567), .C2(net11894), .A(n2871), 
        .ZN(n1145) );
  NOR2_X1 U74 ( .A1(n2530), .A2(n2534), .ZN(n2517) );
  OAI22_X2 U75 ( .A1(n2439), .A2(n54), .B1(n997), .B2(n989), .ZN(n1356) );
  OAI221_X2 U76 ( .B1(n2440), .B2(n3116), .C1(n577), .C2(n50), .A(n612), .ZN(
        n1125) );
  OR2_X4 U77 ( .A1(net11742), .A2(n2616), .ZN(n2621) );
  AOI21_X2 U78 ( .B1(n2441), .B2(net11175), .A(n2446), .ZN(n2442) );
  INV_X4 U79 ( .A(net12968), .ZN(n2441) );
  INV_X2 U80 ( .A(n2442), .ZN(n2606) );
  AOI21_X1 U81 ( .B1(n1073), .B2(n2595), .A(n828), .ZN(n2443) );
  INV_X4 U82 ( .A(n2443), .ZN(goS8) );
  INV_X4 U83 ( .A(net10765), .ZN(n2595) );
  OAI22_X2 U84 ( .A1(n2444), .A2(n54), .B1(n999), .B2(n989), .ZN(n1357) );
  OAI221_X2 U85 ( .B1(n2445), .B2(n3116), .C1(n577), .C2(n49), .A(n606), .ZN(
        n1124) );
  OAI221_X1 U86 ( .B1(n2909), .B2(n2470), .C1(n2908), .C2(net11750), .A(n2907), 
        .ZN(n1135) );
  AOI22_X1 U87 ( .A1(n2638), .A2(U112_DATA1_2), .B1(n2880), .B2(n2639), .ZN(
        n2446) );
  OAI21_X2 U88 ( .B1(n2560), .B2(n2612), .A(n2570), .ZN(n2620) );
  INV_X2 U89 ( .A(n2448), .ZN(n2560) );
  NOR2_X1 U90 ( .A1(n2557), .A2(n2969), .ZN(n2970) );
  OAI22_X2 U91 ( .A1(n2447), .A2(n54), .B1(n995), .B2(n989), .ZN(n1355) );
  NAND3_X1 U92 ( .A1(net10884), .A2(n2520), .A3(n2555), .ZN(n2522) );
  OAI21_X1 U93 ( .B1(net11384), .B2(net11171), .A(U112_DATA1_4), .ZN(n2448) );
  OAI22_X2 U94 ( .A1(n2808), .A2(n2900), .B1(n2603), .B2(n2809), .ZN(n2810) );
  INV_X4 U95 ( .A(n2807), .ZN(n2603) );
  OAI22_X1 U96 ( .A1(net13012), .A2(n181), .B1(n165), .B2(net10761), .ZN(n2775) );
  NAND2_X2 U97 ( .A1(net11403), .A2(U92_DATA2_0), .ZN(n2627) );
  NAND4_X2 U98 ( .A1(n2465), .A2(n2449), .A3(n2461), .A4(n2466), .ZN(n912) );
  OAI211_X2 U99 ( .C1(net11226), .C2(n1020), .A(n2833), .B(r572_A_0_), .ZN(
        n2838) );
  OAI221_X1 U100 ( .B1(n2499), .B2(net11742), .C1(net11121), .C2(net11894), 
        .A(n2918), .ZN(n1131) );
  AOI22_X2 U101 ( .A1(n2635), .A2(U112_DATA1_10), .B1(n2648), .B2(n2908), .ZN(
        n2647) );
  NAND4_X2 U102 ( .A1(n2478), .A2(U91_DATA2_0), .A3(U91_DATA2_1), .A4(n2536), 
        .ZN(n2537) );
  NAND3_X2 U103 ( .A1(n2484), .A2(n2485), .A3(n2524), .ZN(n2548) );
  NAND3_X2 U104 ( .A1(n33), .A2(n2641), .A3(n2813), .ZN(n1068) );
  AOI221_X2 U105 ( .B1(U37_DATA1_0), .B2(n2566), .C1(U37_DATA2_0), .C2(n2473), 
        .A(n2791), .ZN(n2794) );
  NOR2_X1 U106 ( .A1(n2557), .A2(n2960), .ZN(n2961) );
  OR2_X4 U107 ( .A1(n2680), .A2(n2449), .ZN(n2681) );
  XOR2_X2 U108 ( .A(n2642), .B(U92_DATA2_7), .Z(n2601) );
  OAI22_X2 U109 ( .A1(n2450), .A2(n54), .B1(n993), .B2(n989), .ZN(n1354) );
  OAI222_X2 U110 ( .A1(n2451), .A2(n261), .B1(n333), .B2(n3068), .C1(n470), 
        .C2(n2565), .ZN(n1400) );
  INV_X4 U111 ( .A(n2573), .ZN(n2451) );
  NOR3_X1 U112 ( .A1(net12979), .A2(net11119), .A3(net10943), .ZN(n2919) );
  NAND2_X2 U117 ( .A1(net11165), .A2(n2615), .ZN(n2570) );
  OAI22_X1 U122 ( .A1(net13012), .A2(n180), .B1(n164), .B2(net10761), .ZN(
        n2771) );
  OR2_X4 U123 ( .A1(n2587), .A2(n2491), .ZN(n2589) );
  NAND4_X2 U124 ( .A1(U91_DATA2_7), .A2(U92_DATA2_4), .A3(U91_DATA2_4), .A4(
        U91_DATA2_5), .ZN(n2538) );
  AOI21_X2 U125 ( .B1(n2554), .B2(n2529), .A(n2484), .ZN(n2452) );
  INV_X4 U126 ( .A(n2452), .ZN(n2519) );
  AOI21_X2 U127 ( .B1(net10922), .B2(net10923), .A(net17910), .ZN(net10913) );
  NAND4_X2 U128 ( .A1(n2468), .A2(n2453), .A3(n2454), .A4(n2459), .ZN(n913) );
  AND4_X4 U129 ( .A1(n2847), .A2(n2933), .A3(n637), .A4(n2851), .ZN(n2582) );
  OR2_X4 U130 ( .A1(n2677), .A2(n2455), .ZN(n2678) );
  OR2_X4 U131 ( .A1(n2683), .A2(n2456), .ZN(n2684) );
  XOR2_X2 U132 ( .A(n2672), .B(net11466), .Z(n2880) );
  OAI21_X2 U133 ( .B1(n2601), .B2(net11316), .A(n2602), .ZN(n2894) );
  OAI22_X2 U134 ( .A1(n2457), .A2(n54), .B1(n988), .B2(n989), .ZN(n1353) );
  XNOR2_X2 U135 ( .A(net11640), .B(n2669), .ZN(n2689) );
  XOR2_X1 U136 ( .A(net15569), .B(net11417), .Z(n2555) );
  AOI22_X2 U137 ( .A1(U3_U6_DATA4_7), .A2(net17910), .B1(inputSRAM_Addr[7]), 
        .B2(net10847), .ZN(net10844) );
  NOR2_X2 U138 ( .A1(n2458), .A2(n909), .ZN(n2581) );
  INV_X4 U139 ( .A(n2818), .ZN(n2458) );
  OR2_X4 U140 ( .A1(n2675), .A2(n2459), .ZN(n2676) );
  OR2_X4 U141 ( .A1(n2678), .A2(n2460), .ZN(n2679) );
  OR2_X4 U142 ( .A1(n2681), .A2(n2461), .ZN(n2682) );
  OR2_X4 U143 ( .A1(n2684), .A2(n2462), .ZN(n2685) );
  XOR2_X1 U144 ( .A(net12620), .B(U92_DATA2_3), .Z(n2671) );
  XOR2_X1 U145 ( .A(net12590), .B(n2619), .Z(n2617) );
  XNOR2_X1 U146 ( .A(n2799), .B(net12730), .ZN(net11119) );
  OAI221_X2 U147 ( .B1(n2463), .B2(n3116), .C1(n577), .C2(n48), .A(n600), .ZN(
        n1123) );
  OAI21_X1 U148 ( .B1(n416), .B2(net11605), .A(n2691), .ZN(n1285) );
  AOI21_X2 U149 ( .B1(n2810), .B2(n2670), .A(n2568), .ZN(n2646) );
  NOR2_X2 U150 ( .A1(state[4]), .A2(state[0]), .ZN(n2655) );
  XOR2_X2 U151 ( .A(net12566), .B(net11311), .Z(n2483) );
  OR2_X4 U152 ( .A1(n2676), .A2(n2464), .ZN(n2677) );
  OR2_X4 U153 ( .A1(n2679), .A2(n2465), .ZN(n2680) );
  OR2_X4 U154 ( .A1(n2682), .A2(n2466), .ZN(n2683) );
  OR4_X4 U155 ( .A1(net10851), .A2(inputSRAM_Data[0]), .A3(inputSRAM_Data[1]), 
        .A4(inputSRAM_Data[2]), .ZN(n1063) );
  XNOR2_X2 U156 ( .A(net11425), .B(net11334), .ZN(net11121) );
  XNOR2_X2 U157 ( .A(n2662), .B(n3000), .ZN(n3002) );
  NAND2_X2 U158 ( .A1(n41), .A2(n2467), .ZN(sub_387_carry_2_) );
  XNOR2_X2 U159 ( .A(n3063), .B(net10898), .ZN(n257) );
  OR2_X4 U160 ( .A1(n2685), .A2(n2468), .ZN(n2686) );
  OAI222_X2 U161 ( .A1(n2952), .A2(n3084), .B1(n34), .B2(net10887), .C1(
        net10950), .C2(n293), .ZN(n1284) );
  OAI21_X2 U162 ( .B1(n2469), .B2(n3038), .A(n3036), .ZN(n3040) );
  INV_X4 U163 ( .A(n3037), .ZN(n2469) );
  INV_X4 U164 ( .A(net17911), .ZN(net10840) );
  NOR2_X2 U165 ( .A1(n2526), .A2(n2527), .ZN(n2521) );
  NAND2_X2 U166 ( .A1(n2606), .A2(n2607), .ZN(net11384) );
  INV_X4 U167 ( .A(net11119), .ZN(n2524) );
  OAI21_X2 U168 ( .B1(n2528), .B2(n2546), .A(n2553), .ZN(n2552) );
  NOR2_X2 U169 ( .A1(n2500), .A2(U112_DATA1_12), .ZN(n2528) );
  OAI21_X2 U170 ( .B1(net12766), .B2(n2500), .A(n2477), .ZN(n2546) );
  NAND2_X2 U171 ( .A1(n2485), .A2(n2524), .ZN(n2535) );
  NOR2_X2 U172 ( .A1(n2524), .A2(n2485), .ZN(n2525) );
  NOR2_X2 U173 ( .A1(n2481), .A2(n2493), .ZN(n2540) );
  NOR2_X2 U174 ( .A1(n2496), .A2(n2487), .ZN(n2541) );
  NOR2_X2 U175 ( .A1(n2491), .A2(n2495), .ZN(n2536) );
  NAND2_X2 U176 ( .A1(n2793), .A2(n2794), .ZN(net11403) );
  AOI221_X2 U177 ( .B1(U37_DATA5_0), .B2(n2471), .C1(U37_DATA6_0), .C2(n2472), 
        .A(n2792), .ZN(n2793) );
  AOI22_X2 U182 ( .A1(net11454), .A2(U92_DATA2_5), .B1(net12921), .B2(n2673), 
        .ZN(net12590) );
  AOI22_X2 U183 ( .A1(net11316), .A2(U91_DATA2_4), .B1(net11431), .B2(n2644), 
        .ZN(n2643) );
  OAI21_X2 U188 ( .B1(n2517), .B2(n2518), .A(n2519), .ZN(n2516) );
  NAND3_X2 U189 ( .A1(net17910), .A2(net11085), .A3(n2939), .ZN(n3045) );
  INV_X4 U194 ( .A(state[0]), .ZN(net10830) );
  NAND2_X2 U195 ( .A1(n2520), .A2(net10884), .ZN(net11750) );
  NAND2_X2 U200 ( .A1(n2520), .A2(net10884), .ZN(net11894) );
  INV_X4 U201 ( .A(n2640), .ZN(n2952) );
  INV_X4 U206 ( .A(net17910), .ZN(net17911) );
  OAI211_X2 U207 ( .C1(net11742), .C2(n2489), .A(n2522), .B(n2523), .ZN(n1134)
         );
  AOI21_X2 U212 ( .B1(workWrite_Dist[11]), .B2(n2551), .A(net11117), .ZN(n2523) );
  AND3_X4 U213 ( .A1(n2625), .A2(n2624), .A3(n418), .ZN(n2471) );
  AND3_X4 U218 ( .A1(mult_add_378_aco_a_0_), .A2(n2624), .A3(n2625), .ZN(n2472) );
  AND3_X4 U219 ( .A1(mult_add_378_aco_a_0_), .A2(net13049), .A3(n2625), .ZN(
        n2473) );
  NAND2_X2 U220 ( .A1(n2521), .A2(net10850), .ZN(net11113) );
  OR2_X4 U229 ( .A1(U112_DATA1_13), .A2(net11126), .ZN(n2477) );
  AND2_X4 U232 ( .A1(n2545), .A2(n2539), .ZN(n2479) );
  AND2_X4 U233 ( .A1(net12943), .A2(net11131), .ZN(n2500) );
  OAI22_X1 U234 ( .A1(net10919), .A2(net17911), .B1(net10920), .B2(net10921), 
        .ZN(n2501) );
  INV_X4 U235 ( .A(net10941), .ZN(net10936) );
  OAI22_X2 U236 ( .A1(n336), .A2(net10835), .B1(n268), .B2(net10834), .ZN(
        net10941) );
  INV_X4 U237 ( .A(net10847), .ZN(net10834) );
  OAI22_X2 U238 ( .A1(net17911), .A2(net12936), .B1(net10936), .B2(net10937), 
        .ZN(net10930) );
  XOR2_X2 U239 ( .A(net10940), .B(net10936), .Z(n267) );
  NAND3_X2 U240 ( .A1(net10849), .A2(n682), .A3(net10851), .ZN(net10847) );
  NAND2_X1 U241 ( .A1(n1054), .A2(net11236), .ZN(net10849) );
  NAND2_X2 U242 ( .A1(n1054), .A2(net12649), .ZN(n682) );
  NAND2_X2 U243 ( .A1(n1054), .A2(net12639), .ZN(net10851) );
  NAND2_X2 U244 ( .A1(net10847), .A2(inputSRAM_Addr[8]), .ZN(net10839) );
  AOI22_X1 U245 ( .A1(net12938), .A2(net17910), .B1(inputSRAM_Addr[0]), .B2(
        net10847), .ZN(net12936) );
  AND3_X1 U246 ( .A1(state[0]), .A2(state[1]), .A3(net10828), .ZN(net12639) );
  NAND3_X1 U247 ( .A1(net10849), .A2(net10850), .A3(net10851), .ZN(n1041) );
  INV_X2 U248 ( .A(net10922), .ZN(net10919) );
  INV_X4 U249 ( .A(net10923), .ZN(net10920) );
  OAI22_X2 U250 ( .A1(n334), .A2(net17911), .B1(n264), .B2(net10834), .ZN(
        net10923) );
  NOR2_X2 U251 ( .A1(net10840), .A2(net10922), .ZN(net10921) );
  OAI22_X2 U252 ( .A1(net10927), .A2(net17911), .B1(n2502), .B2(n2503), .ZN(
        net10922) );
  INV_X4 U253 ( .A(n2501), .ZN(net10911) );
  INV_X2 U254 ( .A(net10930), .ZN(net10927) );
  INV_X4 U255 ( .A(net10931), .ZN(n2502) );
  OAI22_X2 U256 ( .A1(n335), .A2(net17911), .B1(n266), .B2(net10834), .ZN(
        net10931) );
  NOR2_X2 U257 ( .A1(net10840), .A2(net10930), .ZN(n2503) );
  NOR2_X2 U258 ( .A1(U3_U6_Z_0), .A2(net10840), .ZN(net10937) );
  INV_X4 U259 ( .A(net12936), .ZN(U3_U6_Z_0) );
  INV_X4 U260 ( .A(n2509), .ZN(net10846) );
  AOI22_X2 U261 ( .A1(net10898), .A2(net10840), .B1(net10899), .B2(net17864), 
        .ZN(n2509) );
  NOR2_X2 U262 ( .A1(net10840), .A2(net10846), .ZN(n2504) );
  XOR2_X2 U263 ( .A(net10846), .B(net10840), .Z(net10893) );
  OAI22_X2 U264 ( .A1(net10903), .A2(net17911), .B1(n2505), .B2(n2506), .ZN(
        net10898) );
  OAI22_X1 U265 ( .A1(n331), .A2(net17911), .B1(n258), .B2(net10834), .ZN(
        net10899) );
  OR2_X4 U266 ( .A1(net10840), .A2(net10898), .ZN(net17864) );
  OAI22_X2 U267 ( .A1(n2509), .A2(net17911), .B1(net10844), .B2(n2504), .ZN(
        net10841) );
  INV_X4 U268 ( .A(n2507), .ZN(net10903) );
  INV_X4 U269 ( .A(net10907), .ZN(n2505) );
  OAI22_X2 U270 ( .A1(n332), .A2(net17911), .B1(n260), .B2(net10834), .ZN(
        net10907) );
  NOR2_X2 U271 ( .A1(net10840), .A2(n2507), .ZN(n2506) );
  OAI22_X2 U272 ( .A1(net10911), .A2(net17911), .B1(n2508), .B2(net10913), 
        .ZN(n2507) );
  INV_X4 U273 ( .A(net10915), .ZN(n2508) );
  OAI22_X2 U274 ( .A1(n333), .A2(net17911), .B1(n262), .B2(net10834), .ZN(
        net10915) );
  NAND2_X2 U275 ( .A1(reset), .A2(n1041), .ZN(n1042) );
  XNOR2_X2 U276 ( .A(n2513), .B(n2510), .ZN(n251) );
  XNOR2_X2 U277 ( .A(net17911), .B(n2511), .ZN(n2513) );
  OAI22_X2 U278 ( .A1(net10837), .A2(net17911), .B1(n2512), .B2(net10839), 
        .ZN(n2511) );
  INV_X4 U279 ( .A(net10841), .ZN(net10837) );
  NOR2_X2 U280 ( .A1(net10840), .A2(net10841), .ZN(n2512) );
  NOR2_X2 U281 ( .A1(n252), .A2(net10834), .ZN(n2510) );
  XNOR2_X1 U282 ( .A(net10842), .B(net10841), .ZN(n253) );
  NAND2_X2 U283 ( .A1(n2514), .A2(n2515), .ZN(net12979) );
  INV_X4 U284 ( .A(net10943), .ZN(net10884) );
  INV_X4 U285 ( .A(net11195), .ZN(net11117) );
  INV_X4 U286 ( .A(U91_DATA2_6), .ZN(n2556) );
  INV_X4 U287 ( .A(n637), .ZN(n2526) );
  INV_X4 U288 ( .A(net11226), .ZN(n2527) );
  INV_X4 U289 ( .A(n2525), .ZN(n2529) );
  NAND3_X2 U290 ( .A1(n2531), .A2(n2532), .A3(n2533), .ZN(n2530) );
  NOR2_X2 U291 ( .A1(n2537), .A2(n2538), .ZN(n2539) );
  NAND2_X2 U292 ( .A1(n2541), .A2(n2540), .ZN(n2542) );
  NAND2_X2 U293 ( .A1(U92_DATA2_7), .A2(U92_DATA2_3), .ZN(n2543) );
  NAND2_X2 U294 ( .A1(U92_DATA2_0), .A2(U91_DATA2_6), .ZN(n2544) );
  NOR3_X2 U295 ( .A1(n2542), .A2(n2543), .A3(n2544), .ZN(n2545) );
  NAND2_X2 U296 ( .A1(n2547), .A2(n2484), .ZN(n2534) );
  NAND2_X2 U297 ( .A1(n2483), .A2(n2548), .ZN(n2518) );
  NAND2_X2 U298 ( .A1(n2552), .A2(net11121), .ZN(n2532) );
  NAND2_X2 U299 ( .A1(n2552), .A2(U112_DATA1_14), .ZN(n2531) );
  NAND2_X2 U300 ( .A1(net11126), .A2(U112_DATA1_13), .ZN(n2553) );
  NAND2_X2 U301 ( .A1(n2535), .A2(n2530), .ZN(n2554) );
  INV_X4 U302 ( .A(net12979), .ZN(n2520) );
  INV_X4 U303 ( .A(net11113), .ZN(n2551) );
  NAND2_X2 U304 ( .A1(net11121), .A2(U112_DATA1_14), .ZN(n2533) );
  NAND2_X2 U305 ( .A1(n2525), .A2(n2535), .ZN(n2547) );
  INV_X4 U306 ( .A(n2516), .ZN(n2549) );
  XNOR2_X2 U307 ( .A(net11311), .B(net11309), .ZN(n2550) );
  INV_X4 U308 ( .A(n2555), .ZN(net11136) );
  INV_X4 U309 ( .A(net10835), .ZN(net17910) );
  AND2_X2 U310 ( .A1(n2626), .A2(n418), .ZN(n2561) );
  OR2_X1 U311 ( .A1(n2617), .A2(n2616), .ZN(n2571) );
  INV_X1 U312 ( .A(n2960), .ZN(n2963) );
  OAI22_X1 U313 ( .A1(n13), .A2(n2687), .B1(n339), .B2(n3045), .ZN(n3041) );
  OAI22_X1 U314 ( .A1(n15), .A2(n2687), .B1(n340), .B2(n3045), .ZN(n3027) );
  OAI22_X1 U315 ( .A1(n17), .A2(n2687), .B1(n341), .B2(n3045), .ZN(n3018) );
  OAI22_X1 U316 ( .A1(n19), .A2(n2687), .B1(n342), .B2(n3045), .ZN(n3010) );
  OAI22_X1 U317 ( .A1(n21), .A2(n2687), .B1(n343), .B2(n3045), .ZN(n3005) );
  OAI22_X1 U318 ( .A1(n23), .A2(n2687), .B1(n344), .B2(n3045), .ZN(n2996) );
  OAI22_X1 U319 ( .A1(n25), .A2(n2687), .B1(n345), .B2(n3045), .ZN(n2987) );
  OAI22_X1 U320 ( .A1(n27), .A2(n2687), .B1(n346), .B2(n3045), .ZN(n2978) );
  OAI22_X1 U321 ( .A1(n29), .A2(n2687), .B1(n347), .B2(n3045), .ZN(n2969) );
  OAI22_X1 U322 ( .A1(n31), .A2(n2687), .B1(n348), .B2(n3045), .ZN(n2960) );
  INV_X4 U323 ( .A(n3045), .ZN(n2936) );
  AOI21_X2 U324 ( .B1(net11316), .B2(U91_DATA2_7), .A(n2569), .ZN(net12566) );
  NOR2_X2 U325 ( .A1(net11473), .A2(U92_DATA2_1), .ZN(n2628) );
  OAI21_X2 U326 ( .B1(U91_DATA2_0), .B2(net11316), .A(net12959), .ZN(n2597) );
  NAND2_X2 U327 ( .A1(net11236), .A2(n2559), .ZN(net11226) );
  NAND2_X2 U328 ( .A1(n1073), .A2(net10803), .ZN(net10835) );
  NAND2_X2 U329 ( .A1(net10885), .A2(n3069), .ZN(net10867) );
  NAND2_X1 U330 ( .A1(state[3]), .A2(state[2]), .ZN(n2815) );
  NAND2_X1 U331 ( .A1(n1057), .A2(state[0]), .ZN(n845) );
  INV_X4 U332 ( .A(net11226), .ZN(net10803) );
  OAI221_X2 U333 ( .B1(n981), .B2(net11226), .C1(net11227), .C2(n2851), .A(
        n2850), .ZN(n2937) );
  OAI221_X1 U334 ( .B1(n2470), .B2(n2876), .C1(net11750), .C2(net11186), .A(
        n2875), .ZN(n1144) );
  INV_X4 U335 ( .A(n2600), .ZN(net13039) );
  NAND3_X1 U336 ( .A1(state[2]), .A2(state[3]), .A3(net12639), .ZN(n3093) );
  OAI22_X1 U337 ( .A1(n249), .A2(net10765), .B1(n233), .B2(net10766), .ZN(
        n2623) );
  NAND4_X1 U338 ( .A1(n3096), .A2(state[0]), .A3(net10828), .A4(n575), .ZN(
        n2818) );
  NOR2_X2 U339 ( .A1(n2568), .A2(n2908), .ZN(n2636) );
  AOI221_X1 U340 ( .B1(U38_DATA1_0), .B2(n2566), .C1(U38_DATA2_0), .C2(n2473), 
        .A(n3118), .ZN(n3119) );
  AOI221_X1 U341 ( .B1(U38_DATA1_1), .B2(n2566), .C1(U38_DATA2_1), .C2(n2473), 
        .A(n3123), .ZN(n3124) );
  AOI221_X1 U342 ( .B1(U38_DATA1_2), .B2(n2566), .C1(U38_DATA2_2), .C2(n2473), 
        .A(n3128), .ZN(n3129) );
  AOI221_X1 U343 ( .B1(U38_DATA1_3), .B2(n2566), .C1(U38_DATA2_3), .C2(n2473), 
        .A(n3133), .ZN(n3134) );
  AOI221_X1 U344 ( .B1(U38_DATA1_4), .B2(n2566), .C1(U38_DATA2_4), .C2(n2473), 
        .A(n3138), .ZN(n3139) );
  AOI221_X1 U345 ( .B1(U38_DATA1_5), .B2(n2566), .C1(U38_DATA2_5), .C2(n2473), 
        .A(n3143), .ZN(n3144) );
  AOI221_X1 U346 ( .B1(U38_DATA1_6), .B2(n2566), .C1(U38_DATA2_6), .C2(n2473), 
        .A(n3148), .ZN(n3149) );
  AOI221_X1 U347 ( .B1(U38_DATA1_7), .B2(n2566), .C1(U38_DATA2_7), .C2(n2473), 
        .A(n3153), .ZN(n3154) );
  AOI221_X1 U348 ( .B1(U37_DATA1_6), .B2(n2566), .C1(U37_DATA2_6), .C2(n2473), 
        .A(n2771), .ZN(n2774) );
  AOI221_X1 U349 ( .B1(U37_DATA1_7), .B2(n2566), .C1(U37_DATA2_7), .C2(n2473), 
        .A(n2770), .ZN(net11498) );
  AOI221_X1 U350 ( .B1(U37_DATA1_5), .B2(n2566), .C1(U37_DATA2_5), .C2(n2473), 
        .A(n2775), .ZN(n2778) );
  AOI221_X1 U351 ( .B1(U37_DATA1_3), .B2(n2566), .C1(U37_DATA2_3), .C2(n2473), 
        .A(n2783), .ZN(n2786) );
  AOI221_X1 U352 ( .B1(U37_DATA1_4), .B2(n2566), .C1(U37_DATA2_4), .C2(n2473), 
        .A(n2779), .ZN(n2782) );
  OR2_X2 U353 ( .A1(n2649), .A2(net11131), .ZN(net12766) );
  INV_X4 U354 ( .A(n2646), .ZN(n2648) );
  XNOR2_X1 U355 ( .A(net11387), .B(U92_DATA2_4), .ZN(net12597) );
  NOR2_X2 U356 ( .A1(n2807), .A2(n2899), .ZN(n2808) );
  AND2_X4 U357 ( .A1(net12639), .A2(n2559), .ZN(n2557) );
  AND2_X4 U358 ( .A1(n2577), .A2(n2695), .ZN(n2558) );
  INV_X4 U359 ( .A(net12578), .ZN(net12959) );
  AND2_X4 U360 ( .A1(state[3]), .A2(net11644), .ZN(n2559) );
  XOR2_X2 U361 ( .A(n2592), .B(n2574), .Z(n2562) );
  OR2_X4 U362 ( .A1(n2615), .A2(net11165), .ZN(n2563) );
  AND2_X4 U363 ( .A1(net11316), .A2(U91_DATA2_3), .ZN(n2564) );
  AND2_X4 U364 ( .A1(n2836), .A2(n2835), .ZN(n2565) );
  AND3_X4 U365 ( .A1(n2625), .A2(net13049), .A3(n418), .ZN(n2566) );
  XNOR2_X2 U366 ( .A(net11403), .B(U92_DATA2_0), .ZN(n2567) );
  AND2_X4 U367 ( .A1(U112_DATA1_9), .A2(n2562), .ZN(n2568) );
  AOI22_X2 U368 ( .A1(net11316), .A2(U92_DATA2_7), .B1(n2642), .B2(n2674), 
        .ZN(net12578) );
  AND2_X4 U369 ( .A1(net12730), .A2(net12569), .ZN(n2569) );
  OR2_X4 U370 ( .A1(U92_DATA2_4), .A2(net11458), .ZN(n2572) );
  AND3_X4 U371 ( .A1(net10884), .A2(n3068), .A3(net11227), .ZN(n2573) );
  XNOR2_X2 U372 ( .A(net11316), .B(U91_DATA2_1), .ZN(n2574) );
  OR2_X4 U373 ( .A1(net11316), .A2(U91_DATA2_3), .ZN(n2575) );
  OR2_X4 U374 ( .A1(U91_DATA2_1), .A2(net11316), .ZN(n2576) );
  AND3_X4 U375 ( .A1(n2833), .A2(net10850), .A3(n3069), .ZN(n2577) );
  AND2_X4 U376 ( .A1(U37_DATA5_7), .A2(n2471), .ZN(n2578) );
  XNOR2_X2 U377 ( .A(net11316), .B(U91_DATA2_4), .ZN(n2579) );
  AND3_X4 U378 ( .A1(n3084), .A2(net10943), .A3(n2769), .ZN(n2580) );
  AND2_X4 U379 ( .A1(net11636), .A2(n2669), .ZN(n2583) );
  NAND4_X4 U380 ( .A1(n2584), .A2(n2585), .A3(n2586), .A4(net11498), .ZN(
        net11316) );
  NAND2_X2 U381 ( .A1(n2587), .A2(n2588), .ZN(net12724) );
  NAND2_X2 U382 ( .A1(n2589), .A2(n2590), .ZN(net15569) );
  NOR2_X2 U383 ( .A1(net13039), .A2(n227), .ZN(n2591) );
  NAND2_X2 U384 ( .A1(n2592), .A2(n2576), .ZN(n2587) );
  XNOR2_X2 U385 ( .A(net11316), .B(n2495), .ZN(net11417) );
  XNOR2_X2 U386 ( .A(n2593), .B(n2579), .ZN(net11131) );
  MUX2_X2 U387 ( .A(workRead1_DataInput[75]), .B(U91_DATA2_3), .S(net11609), 
        .Z(n1315) );
  NOR2_X2 U388 ( .A1(n2591), .A2(n2578), .ZN(n2584) );
  NOR2_X2 U389 ( .A1(U91_DATA2_1), .A2(U91_DATA2_2), .ZN(n2594) );
  NAND2_X2 U390 ( .A1(U37_DATA6_7), .A2(n2472), .ZN(n2585) );
  NAND2_X2 U391 ( .A1(n2596), .A2(n2595), .ZN(n2586) );
  INV_X4 U392 ( .A(net11316), .ZN(net11312) );
  NAND2_X2 U393 ( .A1(net11316), .A2(U91_DATA2_0), .ZN(n2598) );
  NAND2_X2 U394 ( .A1(n2598), .A2(n2597), .ZN(n2592) );
  NAND2_X2 U395 ( .A1(net11316), .A2(U91_DATA2_1), .ZN(n2588) );
  NAND2_X2 U396 ( .A1(n2594), .A2(n2587), .ZN(n2599) );
  NAND2_X2 U397 ( .A1(n2599), .A2(net11316), .ZN(n2590) );
  INV_X4 U398 ( .A(n2593), .ZN(net11431) );
  INV_X1 U399 ( .A(net10766), .ZN(n2600) );
  INV_X4 U400 ( .A(n2595), .ZN(net11856) );
  NOR2_X2 U401 ( .A1(U112_DATA1_11), .A2(net11136), .ZN(n2650) );
  OAI221_X1 U418 ( .B1(net11742), .B2(n2904), .C1(n2562), .C2(net11750), .A(
        n2903), .ZN(n1136) );
  NAND2_X2 U419 ( .A1(n2810), .A2(n2670), .ZN(n2652) );
  NOR2_X1 U420 ( .A1(net11113), .A2(n2916), .ZN(n2917) );
  NAND3_X1 U421 ( .A1(state[4]), .A2(net10830), .A3(n2656), .ZN(n3092) );
  NAND3_X1 U422 ( .A1(n1057), .A2(reset), .A3(net10830), .ZN(n2826) );
  NAND2_X1 U423 ( .A1(n1057), .A2(net10830), .ZN(n2817) );
  NAND3_X2 U424 ( .A1(state[1]), .A2(net10828), .A3(net10830), .ZN(net11623)
         );
  NAND2_X2 U425 ( .A1(n2601), .A2(net11316), .ZN(n2602) );
  INV_X4 U426 ( .A(n2617), .ZN(n2622) );
  OAI22_X1 U429 ( .A1(n182), .A2(net13012), .B1(n166), .B2(net10761), .ZN(
        n2779) );
  OAI22_X1 U430 ( .A1(n183), .A2(net13012), .B1(n167), .B2(net10761), .ZN(
        n2783) );
  OAI22_X1 U431 ( .A1(n184), .A2(net10760), .B1(n168), .B2(net10761), .ZN(
        n2787) );
  BUF_X4 U432 ( .A(n416), .Z(net13049) );
  INV_X2 U433 ( .A(n416), .ZN(n2624) );
  OAI221_X1 U434 ( .B1(n2470), .B2(n2486), .C1(net11894), .C2(net11126), .A(
        n2915), .ZN(n1132) );
  NAND2_X2 U435 ( .A1(n2652), .A2(n2636), .ZN(n2635) );
  NAND3_X1 U436 ( .A1(n1054), .A2(state[1]), .A3(state[4]), .ZN(n1040) );
  NAND4_X1 U437 ( .A1(state[4]), .A2(n1054), .A3(state[1]), .A4(state[0]), 
        .ZN(n844) );
  AOI22_X2 U438 ( .A1(n3005), .A2(n2557), .B1(n3000), .B2(n2605), .ZN(n2604)
         );
  OR2_X4 U439 ( .A1(n2557), .A2(n3005), .ZN(n2605) );
  NOR2_X1 U440 ( .A1(net11623), .A2(n2815), .ZN(n2692) );
  NOR3_X1 U441 ( .A1(n828), .A2(net11226), .A3(net13049), .ZN(net11631) );
  NAND2_X1 U442 ( .A1(n2582), .A2(net11226), .ZN(n2848) );
  OAI22_X2 U443 ( .A1(net11375), .A2(n2493), .B1(net12590), .B2(n2797), .ZN(
        n2642) );
  NAND2_X2 U444 ( .A1(n2608), .A2(n2609), .ZN(net12921) );
  NAND2_X2 U445 ( .A1(n2610), .A2(n2611), .ZN(net11368) );
  NOR2_X2 U446 ( .A1(n2613), .A2(n2614), .ZN(n2612) );
  XNOR2_X2 U447 ( .A(net12597), .B(net11458), .ZN(n2614) );
  MUX2_X2 U448 ( .A(U112_DATA1_6), .B(workRead2_DataInput[70]), .S(net11754), 
        .Z(n307) );
  NAND2_X2 U449 ( .A1(net11387), .A2(n2572), .ZN(n2609) );
  NAND2_X2 U450 ( .A1(net11458), .A2(U92_DATA2_4), .ZN(n2608) );
  NAND2_X2 U451 ( .A1(net12968), .A2(U112_DATA1_3), .ZN(n2607) );
  NAND3_X2 U452 ( .A1(n2563), .A2(n2571), .A3(n2620), .ZN(n2611) );
  NAND2_X2 U453 ( .A1(n2617), .A2(n2616), .ZN(n2610) );
  INV_X4 U454 ( .A(n2615), .ZN(net12722) );
  INV_X4 U455 ( .A(n2614), .ZN(net11171) );
  XNOR2_X2 U456 ( .A(U92_DATA2_5), .B(net11454), .ZN(n2618) );
  XNOR2_X2 U457 ( .A(net11450), .B(U92_DATA2_6), .ZN(n2619) );
  XNOR2_X1 U458 ( .A(n2618), .B(net12921), .ZN(n2615) );
  OAI211_X2 U459 ( .C1(n2622), .C2(net11894), .A(n2621), .B(net11162), .ZN(
        n1139) );
  INV_X1 U460 ( .A(net11384), .ZN(n2613) );
  AOI221_X2 U461 ( .B1(U37_DATA5_1), .B2(n2471), .C1(U37_DATA6_1), .C2(n2472), 
        .A(n2623), .ZN(net11475) );
  NAND2_X2 U462 ( .A1(net11475), .A2(net11474), .ZN(net11473) );
  NAND2_X2 U463 ( .A1(n2482), .A2(mult_add_378_aco_a_2_), .ZN(net10765) );
  NAND2_X2 U464 ( .A1(n2482), .A2(net13049), .ZN(net10760) );
  INV_X4 U465 ( .A(n417), .ZN(n2626) );
  INV_X1 U466 ( .A(n2626), .ZN(n2625) );
  NAND3_X1 U467 ( .A1(net10803), .A2(net11227), .A3(mult_add_378_aco_a_0_), 
        .ZN(net11640) );
  MUX2_X2 U468 ( .A(net11640), .B(mult_add_378_aco_a_0_), .S(net11632), .Z(
        n1287) );
  OAI22_X2 U469 ( .A1(net11668), .A2(net11581), .B1(n249), .B2(net11700), .ZN(
        n1185) );
  OAI22_X2 U470 ( .A1(net11405), .A2(n2496), .B1(n2628), .B2(n2627), .ZN(
        net13034) );
  INV_X2 U471 ( .A(net11473), .ZN(net11405) );
  XNOR2_X2 U472 ( .A(n2630), .B(net11405), .ZN(net11399) );
  XNOR2_X2 U473 ( .A(net13082), .B(U92_DATA2_1), .ZN(n2630) );
  AOI221_X2 U474 ( .B1(U37_DATA1_1), .B2(n2566), .C1(U37_DATA2_1), .C2(n2473), 
        .A(n2629), .ZN(net11474) );
  OAI22_X2 U475 ( .A1(n185), .A2(net10760), .B1(n169), .B2(net10761), .ZN(
        n2629) );
  NOR2_X2 U476 ( .A1(net11117), .A2(n2631), .ZN(net11162) );
  NOR2_X2 U477 ( .A1(net11113), .A2(net11164), .ZN(n2631) );
  OAI21_X2 U478 ( .B1(n2632), .B2(n2633), .A(n2634), .ZN(net11195) );
  INV_X4 U479 ( .A(net10942), .ZN(n2634) );
  NAND2_X1 U480 ( .A1(n2634), .A2(n929), .ZN(n930) );
  NAND2_X2 U481 ( .A1(n2634), .A2(net10887), .ZN(net10950) );
  NAND2_X2 U482 ( .A1(n2634), .A2(net10867), .ZN(net10881) );
  NAND4_X2 U483 ( .A1(n664), .A2(n665), .A3(n662), .A4(n663), .ZN(n2633) );
  NAND4_X2 U484 ( .A1(n668), .A2(n669), .A3(n666), .A4(n667), .ZN(n2632) );
  NAND2_X2 U485 ( .A1(net11403), .A2(U92_DATA2_0), .ZN(net13082) );
  OAI22_X1 U486 ( .A1(n11), .A2(n2687), .B1(n338), .B2(n3045), .ZN(n3046) );
  OR2_X1 U487 ( .A1(n2639), .A2(n2880), .ZN(n2638) );
  NAND2_X1 U488 ( .A1(net10803), .A2(reset), .ZN(net10943) );
  NAND2_X2 U489 ( .A1(n2561), .A2(mult_add_378_aco_a_2_), .ZN(net10766) );
  OAI22_X2 U490 ( .A1(n2801), .A2(n2476), .B1(net12620), .B2(n2796), .ZN(
        net11387) );
  INV_X1 U491 ( .A(net10760), .ZN(net13011) );
  INV_X4 U492 ( .A(net13011), .ZN(net13012) );
  XNOR2_X1 U493 ( .A(net13034), .B(U92_DATA2_2), .ZN(n2672) );
  NAND2_X2 U494 ( .A1(n2789), .A2(n2637), .ZN(net12622) );
  AND2_X2 U495 ( .A1(n2790), .A2(n2487), .ZN(n2637) );
  INV_X1 U496 ( .A(n2894), .ZN(n2805) );
  NOR2_X2 U497 ( .A1(n2894), .A2(U112_DATA1_7), .ZN(n2804) );
  OAI22_X1 U498 ( .A1(n2876), .A2(net11399), .B1(n2803), .B2(n2802), .ZN(n2639) );
  AOI22_X2 U499 ( .A1(n2641), .A2(n2557), .B1(graphRead2_Addr[0]), .B2(n2936), 
        .ZN(n2640) );
  OAI22_X2 U500 ( .A1(n2489), .A2(n2555), .B1(n2647), .B2(n2650), .ZN(net12943) );
  XOR2_X2 U501 ( .A(net12724), .B(n2645), .Z(n2908) );
  OAI221_X1 U502 ( .B1(n2470), .B2(n2881), .C1(n2880), .C2(net11750), .A(n2879), .ZN(n1143) );
  OR2_X4 U504 ( .A1(U91_DATA2_4), .A2(net11316), .ZN(n2644) );
  OAI22_X1 U505 ( .A1(n246), .A2(net11856), .B1(n230), .B2(net13039), .ZN(
        n2780) );
  AOI221_X1 U508 ( .B1(U37_DATA5_3), .B2(n2471), .C1(U37_DATA6_3), .C2(n2472), 
        .A(n2784), .ZN(n2785) );
  XNOR2_X2 U509 ( .A(net11316), .B(U91_DATA2_2), .ZN(n2645) );
  OAI22_X1 U510 ( .A1(n245), .A2(net11856), .B1(n229), .B2(net13039), .ZN(
        n2776) );
  OAI22_X1 U511 ( .A1(n248), .A2(net11856), .B1(n232), .B2(net13039), .ZN(
        n2788) );
  OAI22_X1 U512 ( .A1(n247), .A2(net11856), .B1(n231), .B2(net13039), .ZN(
        n2784) );
  OAI22_X1 U513 ( .A1(n244), .A2(net11856), .B1(n228), .B2(net13039), .ZN(
        n2772) );
  AND3_X1 U514 ( .A1(n575), .A2(state[0]), .A3(net10828), .ZN(net12649) );
  AND2_X4 U515 ( .A1(net10803), .A2(n3116), .ZN(n2653) );
  NAND2_X1 U516 ( .A1(net10840), .A2(n2595), .ZN(n2695) );
  XOR2_X1 U517 ( .A(n2661), .B(n2604), .Z(n3007) );
  XOR2_X1 U518 ( .A(n2663), .B(n2998), .Z(n2993) );
  XOR2_X1 U519 ( .A(n2664), .B(n2989), .Z(n2984) );
  XOR2_X1 U520 ( .A(n2667), .B(n2962), .Z(n2957) );
  XOR2_X1 U521 ( .A(n2960), .B(n2687), .Z(n2667) );
  AND3_X1 U522 ( .A1(net10803), .A2(mult_add_378_aco_a_1_), .A3(net11227), 
        .ZN(n2669) );
  XNOR2_X2 U523 ( .A(n2671), .B(n2801), .ZN(net12968) );
  OR2_X1 U524 ( .A1(U92_DATA2_5), .A2(net11454), .ZN(n2673) );
  OAI22_X2 U525 ( .A1(net11312), .A2(n2556), .B1(net11335), .B2(n2651), .ZN(
        net12730) );
  NOR2_X1 U526 ( .A1(U91_DATA2_6), .A2(net11316), .ZN(n2651) );
  AOI221_X2 U527 ( .B1(graphRead1_Addr[7]), .B2(net10863), .C1(U8_DATA3_7), 
        .C2(n3086), .A(n3078), .ZN(n3079) );
  AOI221_X2 U528 ( .B1(graphRead1_Addr[6]), .B2(net10863), .C1(U8_DATA3_6), 
        .C2(n3086), .A(n3076), .ZN(n3077) );
  AOI221_X2 U529 ( .B1(graphRead1_Addr[5]), .B2(net10863), .C1(U8_DATA3_5), 
        .C2(n3086), .A(n3080), .ZN(n3081) );
  AOI221_X2 U530 ( .B1(graphRead1_Addr[4]), .B2(net10863), .C1(U8_DATA3_4), 
        .C2(n3086), .A(n3082), .ZN(n3083) );
  AOI221_X2 U531 ( .B1(graphRead1_Addr[3]), .B2(net10863), .C1(U8_DATA3_3), 
        .C2(n3086), .A(n3085), .ZN(n3087) );
  AOI221_X2 U532 ( .B1(graphRead1_Addr[2]), .B2(net10863), .C1(U8_DATA3_2), 
        .C2(n3086), .A(n3074), .ZN(n3075) );
  AOI221_X2 U533 ( .B1(graphRead1_Addr[1]), .B2(net10863), .C1(U8_DATA3_1), 
        .C2(n3086), .A(n3072), .ZN(n3073) );
  MUX2_X1 U534 ( .A(U112_DATA1_3), .B(workRead2_DataInput[67]), .S(net11754), 
        .Z(n310) );
  NAND4_X1 U535 ( .A1(n1040), .A2(output_WE), .A3(n3092), .A4(n3091), .ZN(
        n1050) );
  XOR2_X1 U537 ( .A(n2658), .B(n3043), .Z(n3033) );
  XOR2_X1 U538 ( .A(n2659), .B(n3020), .Z(n3015) );
  XOR2_X1 U539 ( .A(n2660), .B(n3029), .Z(n3024) );
  XOR2_X1 U540 ( .A(n2665), .B(n2980), .Z(n2975) );
  XOR2_X1 U541 ( .A(n2666), .B(n2971), .Z(n2966) );
  OAI22_X2 U542 ( .A1(n2489), .A2(n2555), .B1(n2647), .B2(n2650), .ZN(n2649)
         );
  OAI221_X1 U543 ( .B1(n277), .B2(net10950), .C1(n19), .C2(net10887), .A(n3006), .ZN(n1276) );
  OAI221_X1 U584 ( .B1(n279), .B2(net10950), .C1(n21), .C2(net10887), .A(n3001), .ZN(n1277) );
  OAI221_X1 U585 ( .B1(n281), .B2(net10950), .C1(n23), .C2(net10887), .A(n2992), .ZN(n1278) );
  OAI221_X1 U586 ( .B1(n283), .B2(net10950), .C1(n25), .C2(net10887), .A(n2983), .ZN(n1279) );
  OAI221_X1 U587 ( .B1(n285), .B2(net10950), .C1(n27), .C2(net10887), .A(n2974), .ZN(n1280) );
  OAI221_X1 U588 ( .B1(n287), .B2(net10950), .C1(n29), .C2(net10887), .A(n2965), .ZN(n1281) );
  OAI221_X1 U589 ( .B1(n289), .B2(net10950), .C1(n31), .C2(net10887), .A(n2956), .ZN(n1282) );
  OAI221_X1 U590 ( .B1(n291), .B2(net10950), .C1(n33), .C2(net10887), .A(n2946), .ZN(n1283) );
  MUX2_X2 U591 ( .A(n3071), .B(net10867), .S(sub_387_A_0_), .Z(n3070) );
  OAI22_X1 U592 ( .A1(n179), .A2(net13012), .B1(n163), .B2(net10761), .ZN(
        n2770) );
  OAI22_X1 U593 ( .A1(n80), .A2(n3084), .B1(n35), .B2(net10867), .ZN(n3078) );
  OAI22_X1 U594 ( .A1(n81), .A2(n3084), .B1(n36), .B2(net10867), .ZN(n3076) );
  OAI22_X1 U595 ( .A1(n82), .A2(n3084), .B1(n37), .B2(net10867), .ZN(n3080) );
  OAI22_X1 U596 ( .A1(n85), .A2(n3084), .B1(n40), .B2(net10867), .ZN(n3074) );
  OAI22_X1 U598 ( .A1(n86), .A2(n3084), .B1(n41), .B2(net10867), .ZN(n3072) );
  OAI22_X1 U599 ( .A1(n83), .A2(n3084), .B1(n38), .B2(net10867), .ZN(n3082) );
  OAI22_X1 U600 ( .A1(n84), .A2(n3084), .B1(n39), .B2(net10867), .ZN(n3085) );
  OAI22_X1 U601 ( .A1(n491), .A2(net10805), .B1(n163), .B2(net11694), .ZN(
        n1255) );
  OAI22_X1 U602 ( .A1(n492), .A2(net10805), .B1(n164), .B2(net11700), .ZN(
        n1254) );
  OAI22_X1 U603 ( .A1(n507), .A2(net10805), .B1(n179), .B2(net11700), .ZN(
        n1239) );
  OAI22_X1 U604 ( .A1(n508), .A2(net10805), .B1(n180), .B2(net11694), .ZN(
        n1238) );
  OAI22_X1 U605 ( .A1(n539), .A2(net10805), .B1(n227), .B2(net11700), .ZN(
        n1207) );
  OAI22_X1 U606 ( .A1(n540), .A2(net10805), .B1(n228), .B2(net11694), .ZN(
        n1206) );
  OAI22_X1 U607 ( .A1(n555), .A2(net10805), .B1(n243), .B2(net11700), .ZN(
        n1191) );
  OAI22_X1 U608 ( .A1(n556), .A2(net10805), .B1(n244), .B2(net11694), .ZN(
        n1190) );
  OAI22_X1 U609 ( .A1(n929), .A2(n87), .B1(n293), .B2(n930), .ZN(n1342) );
  OAI22_X1 U610 ( .A1(n929), .A2(n80), .B1(n279), .B2(n930), .ZN(n1335) );
  OAI22_X1 U611 ( .A1(n929), .A2(n81), .B1(n281), .B2(n930), .ZN(n1336) );
  OAI22_X1 U612 ( .A1(n929), .A2(n82), .B1(n283), .B2(n930), .ZN(n1337) );
  OAI22_X1 U613 ( .A1(n929), .A2(n83), .B1(n285), .B2(n930), .ZN(n1338) );
  OAI22_X1 U614 ( .A1(n929), .A2(n84), .B1(n287), .B2(n930), .ZN(n1339) );
  OAI22_X1 U615 ( .A1(n929), .A2(n85), .B1(n289), .B2(n930), .ZN(n1340) );
  OAI22_X1 U616 ( .A1(n929), .A2(n86), .B1(n291), .B2(n930), .ZN(n1341) );
  OR2_X1 U617 ( .A1(n2562), .A2(U112_DATA1_9), .ZN(n2670) );
  INV_X4 U620 ( .A(net10805), .ZN(net11682) );
  INV_X4 U621 ( .A(n425), .ZN(n3159) );
  INV_X4 U622 ( .A(n2558), .ZN(net11700) );
  INV_X4 U623 ( .A(n2558), .ZN(net11696) );
  INV_X4 U624 ( .A(n2558), .ZN(net11694) );
  INV_X4 U627 ( .A(n2557), .ZN(n2687) );
  INV_X4 U628 ( .A(n849), .ZN(net11609) );
  INV_X4 U629 ( .A(net11516), .ZN(net11754) );
  INV_X4 U630 ( .A(n3084), .ZN(n3049) );
  NAND2_X1 U631 ( .A1(n2845), .A2(net11226), .ZN(n3115) );
  NAND2_X2 U633 ( .A1(n3093), .A2(n3159), .ZN(n424) );
  NAND2_X2 U634 ( .A1(n2694), .A2(net11516), .ZN(n849) );
  OAI21_X2 U635 ( .B1(n563), .B2(n2692), .A(reset), .ZN(n2694) );
  AND2_X1 U636 ( .A1(n2848), .A2(reset), .ZN(n2654) );
  NAND2_X2 U637 ( .A1(n2819), .A2(reset), .ZN(n830) );
  NAND2_X2 U638 ( .A1(n2557), .A2(reset), .ZN(n3084) );
  NAND2_X1 U639 ( .A1(reset), .A2(net10849), .ZN(n1058) );
  OAI211_X1 U640 ( .C1(n1022), .C2(net11226), .A(net10850), .B(n2668), .ZN(
        n3095) );
  NAND2_X2 U641 ( .A1(n2938), .A2(n3045), .ZN(n3053) );
  NAND3_X2 U642 ( .A1(n3036), .A2(reset), .A3(n2935), .ZN(n3038) );
  AND2_X1 U643 ( .A1(n1011), .A2(n575), .ZN(n2656) );
  NAND4_X1 U644 ( .A1(n3096), .A2(net10828), .A3(n575), .A4(net10830), .ZN(
        n3113) );
  XNOR2_X2 U645 ( .A(n3048), .B(n3047), .ZN(n2657) );
  OAI21_X2 U646 ( .B1(n932), .B2(n931), .A(net10850), .ZN(n929) );
  XOR2_X2 U647 ( .A(n3041), .B(n2687), .Z(n2658) );
  XOR2_X2 U648 ( .A(n3018), .B(n2687), .Z(n2659) );
  XOR2_X2 U649 ( .A(n3027), .B(n2687), .Z(n2660) );
  XOR2_X2 U651 ( .A(n3010), .B(n2687), .Z(n2661) );
  XOR2_X2 U652 ( .A(n3005), .B(n2687), .Z(n2662) );
  INV_X4 U653 ( .A(reset), .ZN(net11648) );
  XOR2_X2 U654 ( .A(n2996), .B(n2687), .Z(n2663) );
  XOR2_X2 U657 ( .A(n2987), .B(n2687), .Z(n2664) );
  XOR2_X2 U661 ( .A(n2978), .B(n2687), .Z(n2665) );
  XOR2_X2 U662 ( .A(n2969), .B(n2687), .Z(n2666) );
  INV_X4 U664 ( .A(n907), .ZN(n364) );
  AND2_X1 U665 ( .A1(n2834), .A2(n2924), .ZN(n2668) );
  OR2_X4 U668 ( .A1(U92_DATA2_7), .A2(net11316), .ZN(n2674) );
  OR2_X4 U669 ( .A1(U91_DATA2_7), .A2(net11316), .ZN(net12569) );
  OAI211_X1 U671 ( .C1(n577), .C2(n47), .A(n594), .B(n595), .ZN(n1122) );
  OAI211_X1 U672 ( .C1(n577), .C2(n43), .A(n578), .B(n579), .ZN(n1121) );
  OAI21_X2 U674 ( .B1(n1005), .B2(n989), .A(n1006), .ZN(n1360) );
  OAI21_X1 U676 ( .B1(n1023), .B2(net11226), .A(n2840), .ZN(n1377) );
  AOI22_X2 U678 ( .A1(n1026), .A2(n1020), .B1(n1021), .B2(n3160), .ZN(n1023)
         );
  OAI21_X1 U680 ( .B1(n1013), .B2(net11226), .A(n2843), .ZN(n1376) );
  AOI22_X2 U682 ( .A1(n1017), .A2(n57), .B1(n1018), .B2(n1019), .ZN(n1013) );
  AOI22_X1 U684 ( .A1(n3159), .A2(outputWrite_Addr[3]), .B1(n364), .B2(
        U16_DATA2_3), .ZN(n904) );
  AOI22_X1 U686 ( .A1(n3159), .A2(outputWrite_Addr[11]), .B1(n364), .B2(
        U16_DATA2_11), .ZN(n896) );
  AOI22_X1 U688 ( .A1(n3159), .A2(outputWrite_Addr[5]), .B1(n364), .B2(
        U16_DATA2_5), .ZN(n902) );
  AOI22_X1 U689 ( .A1(n3159), .A2(outputWrite_Addr[10]), .B1(n364), .B2(
        U16_DATA2_10), .ZN(n897) );
  AOI22_X1 U690 ( .A1(n3159), .A2(outputWrite_Addr[4]), .B1(n364), .B2(
        U16_DATA2_4), .ZN(n903) );
  AOI22_X1 U691 ( .A1(n3159), .A2(outputWrite_Addr[12]), .B1(n364), .B2(
        U16_DATA2_12), .ZN(n895) );
  AOI22_X1 U702 ( .A1(n3159), .A2(outputWrite_Addr[6]), .B1(n364), .B2(
        U16_DATA2_6), .ZN(n901) );
  AOI22_X1 U703 ( .A1(n3159), .A2(outputWrite_Addr[7]), .B1(n364), .B2(
        U16_DATA2_7), .ZN(n900) );
  AOI22_X1 U704 ( .A1(n3159), .A2(outputWrite_Addr[8]), .B1(n364), .B2(
        U16_DATA2_8), .ZN(n899) );
  AOI22_X1 U705 ( .A1(n3159), .A2(outputWrite_Addr[1]), .B1(n364), .B2(
        U16_DATA2_1), .ZN(n906) );
  AOI22_X1 U706 ( .A1(n3159), .A2(outputWrite_Addr[9]), .B1(n364), .B2(
        U16_DATA2_9), .ZN(n898) );
  AOI22_X1 U707 ( .A1(n3159), .A2(outputWrite_Addr[2]), .B1(n364), .B2(
        U16_DATA2_2), .ZN(n905) );
  AOI22_X1 U708 ( .A1(n3159), .A2(outputWrite_Addr[13]), .B1(n364), .B2(
        U16_DATA2_13), .ZN(n893) );
  OAI21_X2 U709 ( .B1(n842), .B2(n2816), .A(reset), .ZN(n831) );
  OAI21_X2 U710 ( .B1(n908), .B2(n909), .A(reset), .ZN(n907) );
  AOI21_X1 U711 ( .B1(n910), .B2(n911), .A(n682), .ZN(n908) );
  OAI21_X2 U712 ( .B1(n2), .B2(n849), .A(n1036), .ZN(n1386) );
  OAI21_X2 U713 ( .B1(n3), .B2(n849), .A(n1035), .ZN(n1385) );
  OAI21_X2 U714 ( .B1(n4), .B2(n849), .A(n1034), .ZN(n1384) );
  OAI21_X2 U715 ( .B1(n5), .B2(n849), .A(n1033), .ZN(n1383) );
  OAI21_X2 U716 ( .B1(n6), .B2(n849), .A(n1032), .ZN(n1382) );
  OAI21_X2 U727 ( .B1(n7), .B2(n849), .A(n1031), .ZN(n1381) );
  OAI21_X2 U728 ( .B1(n8), .B2(n849), .A(n1030), .ZN(n1380) );
  OAI21_X2 U729 ( .B1(n9), .B2(n849), .A(n1029), .ZN(n1379) );
  AOI22_X2 U730 ( .A1(n1061), .A2(reset), .B1(n421), .B2(zeroFlag), .ZN(n1060)
         );
  OAI21_X2 U731 ( .B1(n1062), .B2(n1063), .A(reset), .ZN(n1061) );
  OAI21_X2 U732 ( .B1(n772), .B2(n59), .A(n774), .ZN(n1016) );
  AOI22_X2 U733 ( .A1(n58), .A2(U38_DATA4_2), .B1(n737), .B2(U38_DATA3_2), 
        .ZN(n762) );
  AOI22_X2 U734 ( .A1(n58), .A2(U38_DATA4_1), .B1(n737), .B2(U38_DATA3_1), 
        .ZN(n767) );
  AOI22_X2 U735 ( .A1(n58), .A2(U38_DATA4_0), .B1(n737), .B2(U38_DATA3_0), 
        .ZN(n773) );
  AOI22_X2 U736 ( .A1(n58), .A2(U38_DATA4_7), .B1(n737), .B2(U38_DATA3_7), 
        .ZN(n736) );
  AOI22_X2 U746 ( .A1(n58), .A2(U38_DATA4_6), .B1(n737), .B2(U38_DATA3_6), 
        .ZN(n742) );
  AOI22_X2 U747 ( .A1(n58), .A2(U38_DATA4_5), .B1(n737), .B2(U38_DATA3_5), 
        .ZN(n747) );
  AOI22_X2 U748 ( .A1(n58), .A2(U38_DATA4_4), .B1(n737), .B2(U38_DATA3_4), 
        .ZN(n752) );
  AOI22_X2 U752 ( .A1(n58), .A2(U38_DATA4_3), .B1(n737), .B2(U38_DATA3_3), 
        .ZN(n757) );
  XNOR2_X2 U760 ( .A(outputWrite_Addr[1]), .B(n365), .ZN(U16_DATA2_1) );
  NAND2_X2 U773 ( .A1(outputWrite_Addr[1]), .A2(outputWrite_Addr[0]), .ZN(
        n2675) );
  XNOR2_X2 U774 ( .A(outputWrite_Addr[2]), .B(n2675), .ZN(U16_DATA2_2) );
  XNOR2_X2 U775 ( .A(outputWrite_Addr[3]), .B(n2676), .ZN(U16_DATA2_3) );
  XNOR2_X2 U777 ( .A(outputWrite_Addr[4]), .B(n2677), .ZN(U16_DATA2_4) );
  XNOR2_X2 U778 ( .A(outputWrite_Addr[5]), .B(n2678), .ZN(U16_DATA2_5) );
  XNOR2_X2 U779 ( .A(outputWrite_Addr[6]), .B(n2679), .ZN(U16_DATA2_6) );
  XNOR2_X2 U780 ( .A(outputWrite_Addr[7]), .B(n2680), .ZN(U16_DATA2_7) );
  XNOR2_X2 U781 ( .A(outputWrite_Addr[8]), .B(n2681), .ZN(U16_DATA2_8) );
  XNOR2_X2 U782 ( .A(outputWrite_Addr[9]), .B(n2682), .ZN(U16_DATA2_9) );
  XNOR2_X2 U783 ( .A(outputWrite_Addr[10]), .B(n2683), .ZN(U16_DATA2_10) );
  XNOR2_X2 U784 ( .A(outputWrite_Addr[11]), .B(n2684), .ZN(U16_DATA2_11) );
  XNOR2_X2 U785 ( .A(outputWrite_Addr[12]), .B(n2685), .ZN(U16_DATA2_12) );
  XNOR2_X2 U786 ( .A(outputWrite_Addr[13]), .B(n2686), .ZN(U16_DATA2_13) );
  OAI221_X1 U787 ( .B1(net11742), .B2(net11175), .C1(net11894), .C2(net12968), 
        .A(n2884), .ZN(n1142) );
  OAI221_X1 U789 ( .B1(net11742), .B2(net11165), .C1(net11894), .C2(net12722), 
        .A(n2890), .ZN(n1140) );
  NOR2_X1 U790 ( .A1(net12979), .A2(n2580), .ZN(n2814) );
  OAI221_X1 U791 ( .B1(n2470), .B2(n2895), .C1(net11750), .C2(n2894), .A(n2893), .ZN(n1138) );
  OAI22_X1 U792 ( .A1(n171), .A2(net13012), .B1(n155), .B2(net10761), .ZN(
        n3153) );
  OAI22_X1 U793 ( .A1(n172), .A2(net13012), .B1(n156), .B2(net10761), .ZN(
        n3148) );
  OAI22_X1 U794 ( .A1(n173), .A2(net13012), .B1(n157), .B2(net10761), .ZN(
        n3143) );
  OAI22_X1 U795 ( .A1(n174), .A2(net13012), .B1(n158), .B2(net10761), .ZN(
        n3138) );
  OAI22_X1 U796 ( .A1(n175), .A2(net13012), .B1(n159), .B2(net10761), .ZN(
        n3133) );
  OAI22_X1 U797 ( .A1(n176), .A2(net13012), .B1(n160), .B2(net10761), .ZN(
        n3128) );
  OAI22_X1 U798 ( .A1(n177), .A2(net13012), .B1(n161), .B2(net10761), .ZN(
        n3123) );
  OAI22_X1 U799 ( .A1(n178), .A2(net13012), .B1(n162), .B2(net10761), .ZN(
        n3118) );
  INV_X1 U800 ( .A(net13039), .ZN(net11085) );
  OAI22_X1 U801 ( .A1(n241), .A2(net11856), .B1(n225), .B2(net13039), .ZN(
        n3122) );
  OAI22_X1 U802 ( .A1(n239), .A2(net11856), .B1(n223), .B2(net13039), .ZN(
        n3132) );
  OAI22_X1 U803 ( .A1(n237), .A2(net11856), .B1(n221), .B2(net13039), .ZN(
        n3142) );
  OAI22_X1 U804 ( .A1(n235), .A2(net11856), .B1(n219), .B2(net13039), .ZN(
        n3152) );
  OAI22_X1 U805 ( .A1(n236), .A2(net11856), .B1(n220), .B2(net13039), .ZN(
        n3147) );
  OAI22_X1 U806 ( .A1(n238), .A2(net11856), .B1(n222), .B2(net13039), .ZN(
        n3137) );
  OAI22_X1 U807 ( .A1(n240), .A2(net11856), .B1(n224), .B2(net13039), .ZN(
        n3127) );
  OAI22_X1 U808 ( .A1(n242), .A2(net11856), .B1(n226), .B2(net13039), .ZN(
        n3117) );
  INV_X4 U809 ( .A(state[4]), .ZN(net10828) );
  INV_X4 U810 ( .A(net11623), .ZN(net11236) );
  INV_X4 U811 ( .A(state[2]), .ZN(net11644) );
  INV_X4 U812 ( .A(n828), .ZN(net11227) );
  NAND2_X2 U813 ( .A1(net12639), .A2(n1011), .ZN(n2833) );
  INV_X4 U814 ( .A(n2833), .ZN(n2688) );
  NAND2_X2 U815 ( .A1(n2688), .A2(reset), .ZN(n2835) );
  NAND2_X2 U816 ( .A1(n2835), .A2(net10943), .ZN(net11605) );
  INV_X4 U817 ( .A(net11605), .ZN(net11632) );
  INV_X4 U818 ( .A(net11640), .ZN(net11636) );
  MUX2_X2 U819 ( .A(n2689), .B(mult_add_378_aco_a_1_), .S(net11632), .Z(n1286)
         );
  NAND2_X2 U820 ( .A1(n2583), .A2(net11605), .ZN(n2690) );
  MUX2_X2 U821 ( .A(n2690), .B(n2583), .S(net11631), .Z(n2691) );
  NAND2_X2 U822 ( .A1(net12649), .A2(n2559), .ZN(n2851) );
  NAND2_X2 U823 ( .A1(n2851), .A2(net17911), .ZN(n2693) );
  NAND2_X2 U824 ( .A1(n2693), .A2(reset), .ZN(net11516) );
  MUX2_X2 U825 ( .A(workRead1_DataInput[80]), .B(add_118_A_16_), .S(net11609), 
        .Z(n1320) );
  MUX2_X2 U826 ( .A(workRead1_DataInput[73]), .B(U91_DATA2_1), .S(net11609), 
        .Z(n1313) );
  MUX2_X2 U827 ( .A(workRead1_DataInput[72]), .B(U91_DATA2_0), .S(net11609), 
        .Z(n1312) );
  MUX2_X2 U828 ( .A(workRead1_DataInput[79]), .B(U91_DATA2_7), .S(net11609), 
        .Z(n1319) );
  MUX2_X2 U829 ( .A(workRead1_DataInput[78]), .B(U91_DATA2_6), .S(net11609), 
        .Z(n1318) );
  MUX2_X2 U830 ( .A(workRead1_DataInput[77]), .B(U91_DATA2_5), .S(net11609), 
        .Z(n1317) );
  MUX2_X2 U831 ( .A(workRead1_DataInput[76]), .B(U91_DATA2_4), .S(net11609), 
        .Z(n1316) );
  MUX2_X2 U832 ( .A(workRead1_DataInput[74]), .B(U91_DATA2_2), .S(net11609), 
        .Z(n1314) );
  MUX2_X2 U833 ( .A(workRead1_DataInput[71]), .B(U92_DATA2_7), .S(net11609), 
        .Z(n1311) );
  MUX2_X2 U834 ( .A(workRead1_DataInput[70]), .B(U92_DATA2_6), .S(net11609), 
        .Z(n1310) );
  MUX2_X2 U835 ( .A(workRead1_DataInput[69]), .B(U92_DATA2_5), .S(net11609), 
        .Z(n1309) );
  MUX2_X2 U836 ( .A(workRead1_DataInput[68]), .B(U92_DATA2_4), .S(net11609), 
        .Z(n1308) );
  MUX2_X2 U837 ( .A(workRead1_DataInput[67]), .B(U92_DATA2_3), .S(net11609), 
        .Z(n1307) );
  MUX2_X2 U838 ( .A(workRead1_DataInput[66]), .B(U92_DATA2_2), .S(net11609), 
        .Z(n1306) );
  MUX2_X2 U839 ( .A(workRead1_DataInput[65]), .B(U92_DATA2_1), .S(net11609), 
        .Z(n1305) );
  MUX2_X2 U840 ( .A(workRead1_DataInput[64]), .B(U92_DATA2_0), .S(net11609), 
        .Z(n1304) );
  INV_X4 U841 ( .A(n1047), .ZN(net10850) );
  NAND2_X2 U842 ( .A1(n828), .A2(net10803), .ZN(n3069) );
  NAND2_X2 U843 ( .A1(net11696), .A2(net11605), .ZN(net10805) );
  OAI22_X2 U844 ( .A1(net11668), .A2(n474), .B1(net11694), .B2(n2696), .ZN(
        n137) );
  INV_X4 U845 ( .A(graphRead2_DataInput[96]), .ZN(n2698) );
  OAI22_X2 U846 ( .A1(net11668), .A2(n2698), .B1(net11700), .B2(n2697), .ZN(
        n154) );
  INV_X4 U847 ( .A(graphRead2_DataInput[80]), .ZN(n2699) );
  OAI22_X2 U848 ( .A1(net11670), .A2(n2699), .B1(n170), .B2(net11696), .ZN(
        n1248) );
  INV_X4 U849 ( .A(graphRead2_DataInput[64]), .ZN(n2700) );
  OAI22_X2 U850 ( .A1(net11670), .A2(n2700), .B1(n186), .B2(net11694), .ZN(
        n1232) );
  INV_X4 U851 ( .A(graphRead2_DataInput[48]), .ZN(n2702) );
  OAI22_X2 U852 ( .A1(net11668), .A2(n2702), .B1(net11700), .B2(n2701), .ZN(
        n202) );
  INV_X4 U853 ( .A(graphRead2_DataInput[32]), .ZN(n2704) );
  OAI22_X2 U854 ( .A1(net11668), .A2(n2704), .B1(net11694), .B2(n2703), .ZN(
        n218) );
  INV_X4 U855 ( .A(graphRead2_DataInput[16]), .ZN(n2705) );
  OAI22_X2 U856 ( .A1(net11668), .A2(n2705), .B1(n234), .B2(net11696), .ZN(
        n1200) );
  INV_X4 U857 ( .A(graphRead2_DataInput[0]), .ZN(n2706) );
  OAI22_X2 U858 ( .A1(net11670), .A2(n2706), .B1(n250), .B2(net11696), .ZN(
        n1184) );
  OAI22_X2 U859 ( .A1(net11670), .A2(n473), .B1(net11694), .B2(net11592), .ZN(
        n135) );
  INV_X4 U860 ( .A(graphRead2_DataInput[97]), .ZN(n2707) );
  OAI22_X2 U861 ( .A1(net11668), .A2(n2707), .B1(net11700), .B2(net11590), 
        .ZN(n153) );
  INV_X4 U862 ( .A(graphRead2_DataInput[81]), .ZN(n2708) );
  OAI22_X2 U863 ( .A1(net11668), .A2(n2708), .B1(n169), .B2(net11700), .ZN(
        n1249) );
  INV_X4 U864 ( .A(graphRead2_DataInput[65]), .ZN(n2709) );
  OAI22_X2 U865 ( .A1(net11668), .A2(n2709), .B1(n185), .B2(net11694), .ZN(
        n1233) );
  INV_X4 U866 ( .A(graphRead2_DataInput[49]), .ZN(n2710) );
  OAI22_X2 U867 ( .A1(net11670), .A2(n2710), .B1(net11696), .B2(net11586), 
        .ZN(n201) );
  INV_X4 U869 ( .A(graphRead2_DataInput[33]), .ZN(n2711) );
  OAI22_X2 U870 ( .A1(net11670), .A2(n2711), .B1(net11700), .B2(net11584), 
        .ZN(n217) );
  INV_X4 U874 ( .A(graphRead2_DataInput[17]), .ZN(n2712) );
  OAI22_X2 U875 ( .A1(net11670), .A2(n2712), .B1(n233), .B2(net11700), .ZN(
        n1201) );
  INV_X4 U876 ( .A(graphRead2_DataInput[1]), .ZN(net11581) );
  OAI22_X2 U877 ( .A1(net11668), .A2(n472), .B1(net11694), .B2(n2713), .ZN(
        n133) );
  INV_X4 U878 ( .A(graphRead2_DataInput[98]), .ZN(n2715) );
  OAI22_X2 U879 ( .A1(net11668), .A2(n2715), .B1(net11700), .B2(n2714), .ZN(
        n152) );
  INV_X4 U880 ( .A(graphRead2_DataInput[82]), .ZN(n2716) );
  OAI22_X2 U881 ( .A1(net11668), .A2(n2716), .B1(n168), .B2(net11696), .ZN(
        n1250) );
  INV_X4 U882 ( .A(graphRead2_DataInput[66]), .ZN(n2717) );
  OAI22_X2 U883 ( .A1(net11668), .A2(n2717), .B1(n184), .B2(net11694), .ZN(
        n1234) );
  INV_X4 U884 ( .A(graphRead2_DataInput[50]), .ZN(n2719) );
  OAI22_X2 U885 ( .A1(net11670), .A2(n2719), .B1(net11694), .B2(n2718), .ZN(
        n200) );
  INV_X4 U886 ( .A(graphRead2_DataInput[34]), .ZN(n2721) );
  OAI22_X2 U887 ( .A1(net11670), .A2(n2721), .B1(net11700), .B2(n2720), .ZN(
        n216) );
  INV_X4 U888 ( .A(graphRead2_DataInput[18]), .ZN(n2722) );
  OAI22_X2 U889 ( .A1(net11670), .A2(n2722), .B1(n232), .B2(net11696), .ZN(
        n1202) );
  INV_X4 U890 ( .A(graphRead2_DataInput[2]), .ZN(n2723) );
  OAI22_X2 U891 ( .A1(net11670), .A2(n2723), .B1(n248), .B2(net11700), .ZN(
        n1186) );
  OAI22_X2 U892 ( .A1(net11670), .A2(n471), .B1(net11694), .B2(n2724), .ZN(
        n131) );
  INV_X4 U893 ( .A(graphRead2_DataInput[99]), .ZN(n2726) );
  OAI22_X2 U894 ( .A1(net11670), .A2(n2726), .B1(net11700), .B2(n2725), .ZN(
        n151) );
  INV_X4 U897 ( .A(graphRead2_DataInput[83]), .ZN(n2727) );
  OAI22_X2 U899 ( .A1(net11668), .A2(n2727), .B1(n167), .B2(net11696), .ZN(
        n1251) );
  INV_X4 U900 ( .A(graphRead2_DataInput[67]), .ZN(n2728) );
  OAI22_X2 U901 ( .A1(net11670), .A2(n2728), .B1(n183), .B2(net11694), .ZN(
        n1235) );
  INV_X4 U902 ( .A(graphRead2_DataInput[51]), .ZN(n2730) );
  OAI22_X2 U903 ( .A1(net11668), .A2(n2730), .B1(net11694), .B2(n2729), .ZN(
        n199) );
  INV_X4 U904 ( .A(graphRead2_DataInput[35]), .ZN(n2732) );
  OAI22_X2 U905 ( .A1(net11670), .A2(n2732), .B1(net11700), .B2(n2731), .ZN(
        n215) );
  INV_X4 U906 ( .A(graphRead2_DataInput[19]), .ZN(n2733) );
  OAI22_X2 U907 ( .A1(net11668), .A2(n2733), .B1(n231), .B2(net11696), .ZN(
        n1203) );
  INV_X4 U908 ( .A(graphRead2_DataInput[3]), .ZN(n2734) );
  OAI22_X2 U909 ( .A1(net11668), .A2(n2734), .B1(n247), .B2(net11700), .ZN(
        n1187) );
  OAI22_X2 U910 ( .A1(net11668), .A2(n470), .B1(net11696), .B2(n2735), .ZN(
        n129) );
  INV_X4 U911 ( .A(graphRead2_DataInput[100]), .ZN(n2737) );
  OAI22_X2 U912 ( .A1(net11668), .A2(n2737), .B1(net11694), .B2(n2736), .ZN(
        n150) );
  INV_X4 U913 ( .A(graphRead2_DataInput[84]), .ZN(n2738) );
  OAI22_X2 U914 ( .A1(net11670), .A2(n2738), .B1(n166), .B2(net11694), .ZN(
        n1252) );
  INV_X4 U915 ( .A(graphRead2_DataInput[68]), .ZN(n2739) );
  OAI22_X2 U916 ( .A1(net11670), .A2(n2739), .B1(n182), .B2(net11696), .ZN(
        n1236) );
  INV_X4 U917 ( .A(graphRead2_DataInput[52]), .ZN(n2741) );
  OAI22_X2 U918 ( .A1(net11670), .A2(n2741), .B1(net11694), .B2(n2740), .ZN(
        n198) );
  INV_X4 U919 ( .A(graphRead2_DataInput[36]), .ZN(n2743) );
  OAI22_X2 U920 ( .A1(net11670), .A2(n2743), .B1(net11696), .B2(n2742), .ZN(
        n214) );
  INV_X4 U921 ( .A(graphRead2_DataInput[20]), .ZN(n2744) );
  OAI22_X2 U922 ( .A1(net11668), .A2(n2744), .B1(n230), .B2(net11700), .ZN(
        n1204) );
  INV_X4 U923 ( .A(graphRead2_DataInput[4]), .ZN(n2745) );
  OAI22_X2 U924 ( .A1(net11668), .A2(n2745), .B1(n246), .B2(net11696), .ZN(
        n1188) );
  OAI22_X2 U925 ( .A1(net11670), .A2(n469), .B1(net11700), .B2(n2746), .ZN(
        n127) );
  INV_X4 U926 ( .A(graphRead2_DataInput[101]), .ZN(n2748) );
  OAI22_X2 U927 ( .A1(net11668), .A2(n2748), .B1(net11694), .B2(n2747), .ZN(
        n149) );
  INV_X4 U928 ( .A(graphRead2_DataInput[85]), .ZN(n2749) );
  OAI22_X2 U929 ( .A1(net11670), .A2(n2749), .B1(n165), .B2(net11694), .ZN(
        n1253) );
  INV_X4 U930 ( .A(graphRead2_DataInput[69]), .ZN(n2750) );
  OAI22_X2 U931 ( .A1(net11668), .A2(n2750), .B1(n181), .B2(net11700), .ZN(
        n1237) );
  INV_X4 U932 ( .A(graphRead2_DataInput[53]), .ZN(n2752) );
  OAI22_X2 U933 ( .A1(net11668), .A2(n2752), .B1(net11700), .B2(n2751), .ZN(
        n197) );
  INV_X4 U934 ( .A(graphRead2_DataInput[37]), .ZN(n2754) );
  OAI22_X2 U935 ( .A1(net11668), .A2(n2754), .B1(net11700), .B2(n2753), .ZN(
        n213) );
  INV_X4 U936 ( .A(graphRead2_DataInput[21]), .ZN(n2755) );
  OAI22_X2 U937 ( .A1(net11670), .A2(n2755), .B1(n229), .B2(net11694), .ZN(
        n1205) );
  INV_X4 U938 ( .A(graphRead2_DataInput[5]), .ZN(n2756) );
  OAI22_X2 U939 ( .A1(net11670), .A2(n2756), .B1(n245), .B2(net11696), .ZN(
        n1189) );
  OAI22_X2 U940 ( .A1(net11668), .A2(n468), .B1(net11694), .B2(n2757), .ZN(
        n125) );
  INV_X4 U941 ( .A(graphRead2_DataInput[102]), .ZN(n2759) );
  OAI22_X2 U942 ( .A1(net11670), .A2(n2759), .B1(net11700), .B2(n2758), .ZN(
        n148) );
  INV_X4 U943 ( .A(graphRead2_DataInput[54]), .ZN(n2761) );
  OAI22_X2 U944 ( .A1(net11668), .A2(n2761), .B1(net11696), .B2(n2760), .ZN(
        n196) );
  INV_X4 U945 ( .A(graphRead2_DataInput[38]), .ZN(n2763) );
  OAI22_X2 U946 ( .A1(net11670), .A2(n2763), .B1(net11696), .B2(n2762), .ZN(
        n212) );
  OAI22_X2 U947 ( .A1(net11670), .A2(n467), .B1(net11694), .B2(n2764), .ZN(
        n112) );
  INV_X4 U948 ( .A(graphRead2_DataInput[103]), .ZN(n2766) );
  OAI22_X2 U949 ( .A1(net11670), .A2(n2766), .B1(net11694), .B2(n2765), .ZN(
        n147) );
  INV_X4 U950 ( .A(graphRead2_DataInput[55]), .ZN(n2767) );
  OAI22_X2 U951 ( .A1(net11668), .A2(n2767), .B1(net11700), .B2(net11520), 
        .ZN(n195) );
  INV_X4 U952 ( .A(graphRead2_DataInput[39]), .ZN(n2768) );
  OAI22_X2 U953 ( .A1(net11670), .A2(n2768), .B1(net11694), .B2(net11518), 
        .ZN(n211) );
  MUX2_X2 U954 ( .A(U112_DATA1_16), .B(workRead2_DataInput[80]), .S(net11754), 
        .Z(n297) );
  MUX2_X2 U955 ( .A(U112_DATA1_15), .B(workRead2_DataInput[79]), .S(net11754), 
        .Z(n298) );
  MUX2_X2 U956 ( .A(U112_DATA1_14), .B(workRead2_DataInput[78]), .S(net11754), 
        .Z(n299) );
  MUX2_X2 U957 ( .A(U112_DATA1_13), .B(workRead2_DataInput[77]), .S(net11754), 
        .Z(n300) );
  MUX2_X2 U958 ( .A(U112_DATA1_12), .B(workRead2_DataInput[76]), .S(net11754), 
        .Z(n301) );
  MUX2_X2 U959 ( .A(U112_DATA1_11), .B(workRead2_DataInput[75]), .S(net11754), 
        .Z(n302) );
  MUX2_X2 U960 ( .A(U112_DATA1_10), .B(workRead2_DataInput[74]), .S(net11754), 
        .Z(n303) );
  MUX2_X2 U961 ( .A(U112_DATA1_9), .B(workRead2_DataInput[73]), .S(net11754), 
        .Z(n304) );
  MUX2_X2 U962 ( .A(U112_DATA1_8), .B(workRead2_DataInput[72]), .S(net11754), 
        .Z(n305) );
  MUX2_X2 U963 ( .A(U112_DATA1_7), .B(workRead2_DataInput[71]), .S(net11754), 
        .Z(n306) );
  MUX2_X2 U964 ( .A(U112_DATA1_5), .B(workRead2_DataInput[69]), .S(net11754), 
        .Z(n308) );
  MUX2_X2 U965 ( .A(U112_DATA1_4), .B(workRead2_DataInput[68]), .S(net11754), 
        .Z(n309) );
  MUX2_X2 U966 ( .A(U112_DATA1_2), .B(workRead2_DataInput[66]), .S(net11754), 
        .Z(n311) );
  MUX2_X2 U967 ( .A(U112_DATA1_0), .B(workRead2_DataInput[64]), .S(net11754), 
        .Z(n313) );
  MUX2_X2 U968 ( .A(U112_DATA1_1), .B(workRead2_DataInput[65]), .S(net11754), 
        .Z(n312) );
  INV_X4 U969 ( .A(n682), .ZN(net11292) );
  NAND2_X2 U970 ( .A1(net11292), .A2(reset), .ZN(n2769) );
  XOR2_X2 U971 ( .A(net11316), .B(U91_DATA2_7), .Z(n2799) );
  AOI221_X2 U972 ( .B1(U37_DATA5_6), .B2(n2471), .C1(U37_DATA6_6), .C2(n2472), 
        .A(n2772), .ZN(n2773) );
  NAND2_X2 U973 ( .A1(n2774), .A2(n2773), .ZN(net11450) );
  INV_X4 U974 ( .A(net11450), .ZN(net11375) );
  AOI221_X2 U975 ( .B1(U37_DATA5_5), .B2(n2471), .C1(U37_DATA6_5), .C2(n2472), 
        .A(n2776), .ZN(n2777) );
  NAND2_X2 U976 ( .A1(n2778), .A2(n2777), .ZN(net11454) );
  AOI221_X2 U977 ( .B1(U37_DATA5_4), .B2(n2471), .C1(U37_DATA6_4), .C2(n2472), 
        .A(n2780), .ZN(n2781) );
  NAND2_X2 U978 ( .A1(n2782), .A2(n2781), .ZN(net11458) );
  NAND2_X2 U979 ( .A1(n2786), .A2(n2785), .ZN(n2795) );
  INV_X4 U980 ( .A(n2795), .ZN(n2801) );
  AOI221_X2 U981 ( .B1(U37_DATA1_2), .B2(n2566), .C1(U37_DATA2_2), .C2(n2473), 
        .A(n2787), .ZN(n2790) );
  AOI221_X2 U982 ( .B1(U37_DATA5_2), .B2(n2471), .C1(U37_DATA6_2), .C2(n2472), 
        .A(n2788), .ZN(n2789) );
  NAND2_X2 U983 ( .A1(n2789), .A2(n2790), .ZN(net11466) );
  OAI22_X2 U984 ( .A1(n186), .A2(net10760), .B1(n170), .B2(net10761), .ZN(
        n2791) );
  OAI22_X2 U985 ( .A1(n250), .A2(net10765), .B1(n234), .B2(net10766), .ZN(
        n2792) );
  NOR2_X2 U986 ( .A1(U92_DATA2_3), .A2(n2795), .ZN(n2796) );
  NOR2_X2 U987 ( .A1(U92_DATA2_6), .A2(net11450), .ZN(n2797) );
  NOR2_X2 U988 ( .A1(U91_DATA2_5), .A2(net11316), .ZN(n2798) );
  OAI22_X2 U989 ( .A1(net11312), .A2(n2497), .B1(n2643), .B2(n2798), .ZN(
        net11425) );
  INV_X4 U990 ( .A(net11425), .ZN(net11335) );
  XOR2_X2 U991 ( .A(net11316), .B(U91_DATA2_5), .Z(n2800) );
  XOR2_X2 U992 ( .A(n2800), .B(n2643), .Z(net11126) );
  INV_X4 U993 ( .A(net11399), .ZN(net11186) );
  NOR2_X2 U994 ( .A1(U112_DATA1_1), .A2(net11186), .ZN(n2803) );
  NAND2_X2 U995 ( .A1(U112_DATA1_0), .A2(n2567), .ZN(n2802) );
  OAI22_X2 U996 ( .A1(n2895), .A2(n2805), .B1(net11368), .B2(n2804), .ZN(n2807) );
  XOR2_X2 U997 ( .A(net11316), .B(U91_DATA2_0), .Z(n2806) );
  XOR2_X2 U998 ( .A(n2806), .B(net12578), .Z(n2899) );
  INV_X4 U999 ( .A(n2899), .ZN(n2809) );
  XOR2_X2 U1000 ( .A(net11316), .B(U91_DATA2_6), .Z(net11334) );
  XOR2_X2 U1001 ( .A(net11316), .B(add_118_A_16_), .Z(net11311) );
  NOR2_X2 U1002 ( .A1(add_118_A_16_), .A2(net11316), .ZN(n2811) );
  OAI22_X2 U1003 ( .A1(net11312), .A2(n2478), .B1(net12566), .B2(n2811), .ZN(
        net11309) );
  NOR2_X2 U1004 ( .A1(net11292), .A2(n2557), .ZN(n2812) );
  OAI22_X2 U1005 ( .A1(n2814), .A2(n2813), .B1(n2580), .B2(n2812), .ZN(n1154)
         );
  INV_X4 U1019 ( .A(n2815), .ZN(n3096) );
  INV_X4 U1020 ( .A(n2818), .ZN(n2816) );
  NAND3_X2 U1021 ( .A1(n845), .A2(n844), .A3(n2817), .ZN(n909) );
  NAND2_X2 U1023 ( .A1(n2581), .A2(net10850), .ZN(n425) );
  INV_X4 U1024 ( .A(n3093), .ZN(n2819) );
  INV_X4 U1025 ( .A(n830), .ZN(n2828) );
  OAI221_X2 U1026 ( .B1(n381), .B2(n424), .C1(n3098), .C2(n2826), .A(n831), 
        .ZN(n2820) );
  AOI221_X2 U1027 ( .B1(n2828), .B2(U92_DATA2_0), .C1(n834), .C2(U97_DATA4_0), 
        .A(n2820), .ZN(n2821) );
  INV_X4 U1028 ( .A(n2821), .ZN(n1303) );
  OAI221_X2 U1029 ( .B1(n380), .B2(n424), .C1(n3100), .C2(n2826), .A(n831), 
        .ZN(n2822) );
  AOI221_X2 U1030 ( .B1(n2828), .B2(U92_DATA2_1), .C1(n834), .C2(U97_DATA4_1), 
        .A(n2822), .ZN(n2823) );
  INV_X4 U1036 ( .A(n2823), .ZN(n1302) );
  OAI221_X2 U1037 ( .B1(n379), .B2(n424), .C1(n3102), .C2(n2826), .A(n831), 
        .ZN(n2824) );
  AOI221_X2 U1038 ( .B1(n2828), .B2(U92_DATA2_2), .C1(n834), .C2(U97_DATA4_2), 
        .A(n2824), .ZN(n2825) );
  INV_X4 U1047 ( .A(n2825), .ZN(n1301) );
  NAND2_X2 U1048 ( .A1(n834), .A2(U97_DATA4_3), .ZN(n2830) );
  INV_X4 U1058 ( .A(n2826), .ZN(n3158) );
  NOR2_X2 U1059 ( .A1(n378), .A2(n424), .ZN(n2827) );
  AOI221_X2 U1094 ( .B1(n2828), .B2(U92_DATA2_3), .C1(n3158), .C2(U97_DATA3_3), 
        .A(n2827), .ZN(n2829) );
  NAND3_X2 U1095 ( .A1(n2830), .A2(n831), .A3(n2829), .ZN(n1300) );
  NAND2_X2 U1096 ( .A1(n1011), .A2(net12649), .ZN(n637) );
  NAND2_X2 U1097 ( .A1(n2656), .A2(n2655), .ZN(n2933) );
  NAND3_X2 U1098 ( .A1(n2687), .A2(n2833), .A3(n2933), .ZN(n2832) );
  NAND3_X2 U1099 ( .A1(n575), .A2(n2559), .A3(n2655), .ZN(n2924) );
  NAND2_X2 U1110 ( .A1(n2924), .A2(n2851), .ZN(n2841) );
  INV_X4 U1111 ( .A(n2841), .ZN(n2845) );
  NAND3_X2 U1112 ( .A1(work_WE), .A2(n2551), .A3(n2845), .ZN(n2831) );
  NAND2_X2 U1113 ( .A1(n2526), .A2(reset), .ZN(net10942) );
  OAI221_X2 U1114 ( .B1(n2832), .B2(n2831), .C1(graphData1_Zero_reg), .C2(
        net10942), .A(net10943), .ZN(n1351) );
  NAND3_X2 U1115 ( .A1(n61), .A2(n60), .A3(n59), .ZN(n735) );
  NAND2_X2 U1142 ( .A1(n982), .A2(n337), .ZN(n2939) );
  NAND3_X2 U1143 ( .A1(n1073), .A2(n735), .A3(n2939), .ZN(n1022) );
  INV_X4 U1144 ( .A(n1020), .ZN(n3160) );
  INV_X4 U1145 ( .A(n2851), .ZN(n2928) );
  NAND2_X2 U1146 ( .A1(n2928), .A2(n1073), .ZN(n2834) );
  NAND2_X2 U1147 ( .A1(net10884), .A2(n828), .ZN(n2836) );
  OAI221_X2 U1158 ( .B1(net11648), .B2(n2668), .C1(n1022), .C2(net10943), .A(
        n2565), .ZN(n2837) );
  INV_X4 U1159 ( .A(n2837), .ZN(n55) );
  MUX2_X2 U1160 ( .A(n2838), .B(r572_A_0_), .S(n55), .Z(n1378) );
  NAND2_X2 U1161 ( .A1(n1025), .A2(n2841), .ZN(n2839) );
  MUX2_X2 U1162 ( .A(n2839), .B(n60), .S(n55), .Z(n2840) );
  NAND2_X2 U1163 ( .A1(n1016), .A2(n2841), .ZN(n2842) );
  MUX2_X2 U1166 ( .A(n2842), .B(n59), .S(n55), .Z(n2843) );
  NAND3_X2 U1167 ( .A1(n2577), .A2(net17911), .A3(n2687), .ZN(n3068) );
  NAND2_X2 U1168 ( .A1(n2573), .A2(net12936), .ZN(n2844) );
  OAI221_X2 U1169 ( .B1(n337), .B2(n3068), .C1(n474), .C2(n2565), .A(n2844), 
        .ZN(n1404) );
  NAND3_X2 U1170 ( .A1(n3115), .A2(reset), .A3(n3095), .ZN(n2846) );
  OAI22_X2 U1171 ( .A1(n768), .A2(n2846), .B1(n103), .B2(n3095), .ZN(n1162) );
  OAI22_X2 U1172 ( .A1(n763), .A2(n2846), .B1(n102), .B2(n3095), .ZN(n1161) );
  OAI22_X2 U1173 ( .A1(n758), .A2(n2846), .B1(n101), .B2(n3095), .ZN(n1160) );
  OAI22_X2 U1174 ( .A1(n753), .A2(n2846), .B1(n100), .B2(n3095), .ZN(n1159) );
  OAI22_X2 U1175 ( .A1(n748), .A2(n2846), .B1(n99), .B2(n3095), .ZN(n1158) );
  OAI22_X2 U1177 ( .A1(n743), .A2(n2846), .B1(n98), .B2(n3095), .ZN(n1157) );
  OAI22_X2 U1179 ( .A1(n738), .A2(n2846), .B1(n97), .B2(n3095), .ZN(n1156) );
  OAI22_X2 U1180 ( .A1(n725), .A2(n2846), .B1(n96), .B2(n3095), .ZN(n1155) );
  MUX2_X2 U1181 ( .A(U113_DATA2_0), .B(workRead2_DataInput[0]), .S(net11754), 
        .Z(n321) );
  NAND2_X2 U1182 ( .A1(n1011), .A2(net11236), .ZN(n2847) );
  NAND2_X2 U1183 ( .A1(n2847), .A2(n2933), .ZN(n2849) );
  NOR3_X2 U1184 ( .A1(n2526), .A2(n1047), .A3(n2849), .ZN(n2850) );
  NAND2_X2 U1185 ( .A1(n2654), .A2(n2937), .ZN(n2866) );
  OAI22_X2 U1186 ( .A1(n445), .A2(n2866), .B1(n53), .B2(n2937), .ZN(n1361) );
  MUX2_X2 U1187 ( .A(U97_DATA2_0), .B(n2852), .S(n2565), .Z(n1352) );
  NAND2_X2 U1188 ( .A1(workWrite_Pred[0]), .A2(n2551), .ZN(n2853) );
  MUX2_X2 U1189 ( .A(U113_DATA2_1), .B(workRead2_DataInput[1]), .S(net11754), 
        .Z(n320) );
  OAI22_X2 U1190 ( .A1(n444), .A2(n2866), .B1(n52), .B2(n2937), .ZN(n1363) );
  MUX2_X2 U1191 ( .A(U97_DATA2_1), .B(n2854), .S(n2565), .Z(n1362) );
  NAND2_X2 U1192 ( .A1(workWrite_Pred[1]), .A2(n2551), .ZN(n2855) );
  MUX2_X2 U1196 ( .A(U113_DATA2_2), .B(workRead2_DataInput[2]), .S(net11754), 
        .Z(n319) );
  OAI22_X2 U1197 ( .A1(n443), .A2(n2866), .B1(n51), .B2(n2937), .ZN(n1365) );
  MUX2_X2 U1198 ( .A(U97_DATA2_2), .B(n2856), .S(n2565), .Z(n1364) );
  NAND2_X2 U1199 ( .A1(workWrite_Pred[2]), .A2(n2551), .ZN(n2857) );
  OAI221_X2 U1201 ( .B1(n396), .B2(net11742), .C1(n67), .C2(net11894), .A(
        n2857), .ZN(n1151) );
  MUX2_X2 U1202 ( .A(U113_DATA2_3), .B(workRead2_DataInput[3]), .S(net11754), 
        .Z(n318) );
  OAI22_X2 U1203 ( .A1(n442), .A2(n2866), .B1(n50), .B2(n2937), .ZN(n1367) );
  MUX2_X2 U1204 ( .A(U97_DATA2_3), .B(n2858), .S(n2565), .Z(n1366) );
  NAND2_X2 U1205 ( .A1(workWrite_Pred[3]), .A2(n2551), .ZN(n2859) );
  MUX2_X2 U1206 ( .A(U113_DATA2_4), .B(workRead2_DataInput[4]), .S(net11754), 
        .Z(n317) );
  OAI22_X2 U1207 ( .A1(n441), .A2(n2866), .B1(n49), .B2(n2937), .ZN(n1369) );
  MUX2_X2 U1208 ( .A(U97_DATA2_4), .B(n2860), .S(n2565), .Z(n1368) );
  NAND2_X2 U1209 ( .A1(workWrite_Pred[4]), .A2(n2551), .ZN(n2861) );
  MUX2_X2 U1210 ( .A(U113_DATA2_5), .B(workRead2_DataInput[5]), .S(net11754), 
        .Z(n316) );
  OAI22_X2 U1211 ( .A1(n440), .A2(n2866), .B1(n48), .B2(n2937), .ZN(n1371) );
  MUX2_X2 U1212 ( .A(U97_DATA2_5), .B(n2862), .S(n2565), .Z(n1370) );
  NAND2_X2 U1213 ( .A1(workWrite_Pred[5]), .A2(n2551), .ZN(n2863) );
  OAI221_X2 U1214 ( .B1(n393), .B2(net11742), .C1(n64), .C2(net11894), .A(
        n2863), .ZN(n1148) );
  MUX2_X2 U1215 ( .A(U113_DATA2_6), .B(workRead2_DataInput[6]), .S(net11754), 
        .Z(n315) );
  OAI22_X2 U1216 ( .A1(n439), .A2(n2866), .B1(n47), .B2(n2937), .ZN(n1373) );
  MUX2_X2 U1217 ( .A(U97_DATA2_6), .B(n2864), .S(n2565), .Z(n1372) );
  NAND2_X2 U1218 ( .A1(workWrite_Pred[6]), .A2(n2551), .ZN(n2865) );
  MUX2_X2 U1219 ( .A(U113_DATA2_7), .B(workRead2_DataInput[7]), .S(net11754), 
        .Z(n314) );
  OAI22_X2 U1220 ( .A1(n438), .A2(n2866), .B1(n43), .B2(n2937), .ZN(n1375) );
  MUX2_X2 U1221 ( .A(U97_DATA2_7), .B(n2867), .S(n2565), .Z(n1374) );
  NAND2_X2 U1222 ( .A1(workWrite_Pred[7]), .A2(n2551), .ZN(n2868) );
  OAI221_X2 U1223 ( .B1(n391), .B2(n2470), .C1(n62), .C2(net11894), .A(n2868), 
        .ZN(n1146) );
  NOR2_X2 U1224 ( .A1(net11113), .A2(n2869), .ZN(n2870) );
  NOR2_X2 U1225 ( .A1(net11117), .A2(n2870), .ZN(n2871) );
  NOR2_X2 U1226 ( .A1(net11113), .A2(n2873), .ZN(n2874) );
  NOR2_X2 U1227 ( .A1(net11117), .A2(n2874), .ZN(n2875) );
  NOR2_X2 U1228 ( .A1(net11113), .A2(n2877), .ZN(n2878) );
  NOR2_X2 U1229 ( .A1(net11117), .A2(n2878), .ZN(n2879) );
  NOR2_X2 U1230 ( .A1(net11113), .A2(n2882), .ZN(n2883) );
  NOR2_X2 U1231 ( .A1(net11117), .A2(n2883), .ZN(n2884) );
  NOR2_X2 U1232 ( .A1(net11113), .A2(n2885), .ZN(n2886) );
  NOR2_X2 U1233 ( .A1(net11117), .A2(n2886), .ZN(n2887) );
  OAI221_X2 U1234 ( .B1(net11170), .B2(net11742), .C1(net11750), .C2(net11171), 
        .A(n2887), .ZN(n1141) );
  NOR2_X2 U1235 ( .A1(net11113), .A2(n2888), .ZN(n2889) );
  NOR2_X2 U1236 ( .A1(net11117), .A2(n2889), .ZN(n2890) );
  NOR2_X2 U1237 ( .A1(net11113), .A2(n2891), .ZN(n2892) );
  NOR2_X2 U1238 ( .A1(net11117), .A2(n2892), .ZN(n2893) );
  NOR2_X2 U1239 ( .A1(net11113), .A2(n2896), .ZN(n2897) );
  NOR2_X2 U1240 ( .A1(net11117), .A2(n2897), .ZN(n2898) );
  OAI221_X2 U1241 ( .B1(n2900), .B2(net11742), .C1(n2899), .C2(net11750), .A(
        n2898), .ZN(n1137) );
  NOR2_X2 U1242 ( .A1(net11113), .A2(n2901), .ZN(n2902) );
  NOR2_X2 U1243 ( .A1(net11117), .A2(n2902), .ZN(n2903) );
  NOR2_X2 U1244 ( .A1(net11113), .A2(n2905), .ZN(n2906) );
  NOR2_X2 U1245 ( .A1(net11117), .A2(n2906), .ZN(n2907) );
  NOR2_X2 U1246 ( .A1(net11113), .A2(n2910), .ZN(n2911) );
  NOR2_X2 U1247 ( .A1(net11117), .A2(n2911), .ZN(n2912) );
  OAI221_X2 U1248 ( .B1(n2488), .B2(net11742), .C1(net11131), .C2(net11750), 
        .A(n2912), .ZN(n1133) );
  NOR2_X2 U1249 ( .A1(net11113), .A2(n2913), .ZN(n2914) );
  NOR2_X2 U1250 ( .A1(net11117), .A2(n2914), .ZN(n2915) );
  NOR2_X2 U1251 ( .A1(net11117), .A2(n2917), .ZN(n2918) );
  NOR2_X2 U1252 ( .A1(n2919), .A2(net11117), .ZN(n2920) );
  OAI221_X2 U1253 ( .B1(net11113), .B2(n2921), .C1(net11742), .C2(n2485), .A(
        n2920), .ZN(n1130) );
  NAND2_X2 U1254 ( .A1(workWrite_Dist[16]), .A2(n2551), .ZN(n2922) );
  INV_X4 U1255 ( .A(n2933), .ZN(n2923) );
  NOR4_X2 U1256 ( .A1(n2526), .A2(n2923), .A3(n1047), .A4(n2557), .ZN(n2930)
         );
  INV_X4 U1257 ( .A(n981), .ZN(n2927) );
  INV_X4 U1258 ( .A(n2924), .ZN(n2926) );
  AND4_X2 U1259 ( .A1(n983), .A2(n982), .A3(net10803), .A4(n735), .ZN(n2925)
         );
  AOI221_X2 U1260 ( .B1(n2928), .B2(n2927), .C1(n2926), .C2(n828), .A(n2925), 
        .ZN(n2929) );
  NAND2_X2 U1261 ( .A1(n2930), .A2(n2929), .ZN(n3036) );
  INV_X4 U1262 ( .A(n3115), .ZN(n2934) );
  INV_X4 U1263 ( .A(graphData1_Zero_reg), .ZN(n2931) );
  NAND2_X2 U1264 ( .A1(n2526), .A2(n2931), .ZN(n2932) );
  NAND3_X2 U1265 ( .A1(n2934), .A2(n2933), .A3(n2932), .ZN(n2935) );
  OAI22_X2 U1266 ( .A1(graphRead1_Addr[0]), .A2(n3038), .B1(n293), .B2(n3036), 
        .ZN(n1350) );
  INV_X4 U1267 ( .A(n929), .ZN(net11093) );
  NAND2_X2 U1268 ( .A1(n2936), .A2(reset), .ZN(n2947) );
  INV_X4 U1269 ( .A(n2937), .ZN(n2938) );
  NAND4_X2 U1270 ( .A1(n2582), .A2(n1073), .A3(net11085), .A4(n2939), .ZN(
        n2940) );
  NAND3_X2 U1271 ( .A1(n2654), .A2(n3053), .A3(n2940), .ZN(n3055) );
  INV_X4 U1272 ( .A(n3055), .ZN(n2941) );
  NAND2_X2 U1273 ( .A1(graphRead1_DataInput[0]), .A2(n2941), .ZN(n2942) );
  OAI221_X2 U1274 ( .B1(n2952), .B2(n2947), .C1(n350), .C2(n3053), .A(n2942), 
        .ZN(n1271) );
  INV_X4 U1275 ( .A(U3_U3_DATA6_1), .ZN(n2943) );
  OAI22_X2 U1276 ( .A1(n3038), .A2(n2943), .B1(n291), .B2(n3036), .ZN(n1349)
         );
  XNOR2_X2 U1277 ( .A(n2952), .B(n2687), .ZN(n2945) );
  OAI22_X2 U1278 ( .A1(n33), .A2(n2687), .B1(n349), .B2(n3045), .ZN(n2944) );
  INV_X4 U1279 ( .A(n2944), .ZN(n2954) );
  XNOR2_X2 U1280 ( .A(n2945), .B(n2954), .ZN(n2948) );
  NAND2_X2 U1281 ( .A1(n3049), .A2(n2948), .ZN(n2946) );
  INV_X4 U1282 ( .A(graphRead1_DataInput[1]), .ZN(n2950) );
  INV_X4 U1283 ( .A(n2947), .ZN(n3051) );
  NAND2_X2 U1284 ( .A1(n3051), .A2(n2948), .ZN(n2949) );
  OAI221_X2 U1285 ( .B1(n3055), .B2(n2950), .C1(n349), .C2(n3053), .A(n2949), 
        .ZN(n1270) );
  INV_X4 U1286 ( .A(U3_U3_DATA6_2), .ZN(n2951) );
  OAI22_X2 U1287 ( .A1(n3038), .A2(n2951), .B1(n289), .B2(n3036), .ZN(n1348)
         );
  NOR2_X2 U1288 ( .A1(n2557), .A2(n2952), .ZN(n2953) );
  OAI22_X2 U1289 ( .A1(n2640), .A2(n2687), .B1(n2954), .B2(n2953), .ZN(n2955)
         );
  INV_X4 U1290 ( .A(n2955), .ZN(n2962) );
  NAND2_X2 U1291 ( .A1(n3049), .A2(n2957), .ZN(n2956) );
  NAND2_X2 U1292 ( .A1(n3051), .A2(n2957), .ZN(n2958) );
  OAI221_X2 U1293 ( .B1(n456), .B2(n3055), .C1(n348), .C2(n3053), .A(n2958), 
        .ZN(n1269) );
  INV_X4 U1294 ( .A(U3_U3_DATA6_3), .ZN(n2959) );
  OAI22_X2 U1295 ( .A1(n3038), .A2(n2959), .B1(n287), .B2(n3036), .ZN(n1347)
         );
  OAI22_X2 U1296 ( .A1(n2963), .A2(n2687), .B1(n2962), .B2(n2961), .ZN(n2964)
         );
  INV_X4 U1297 ( .A(n2964), .ZN(n2971) );
  NAND2_X2 U1298 ( .A1(n3049), .A2(n2966), .ZN(n2965) );
  NAND2_X2 U1299 ( .A1(n3051), .A2(n2966), .ZN(n2967) );
  OAI221_X2 U1300 ( .B1(n455), .B2(n3055), .C1(n347), .C2(n3053), .A(n2967), 
        .ZN(n1268) );
  INV_X4 U1301 ( .A(U3_U3_DATA6_4), .ZN(n2968) );
  OAI22_X2 U1302 ( .A1(n3038), .A2(n2968), .B1(n285), .B2(n3036), .ZN(n1346)
         );
  INV_X4 U1303 ( .A(n2969), .ZN(n2972) );
  OAI22_X2 U1304 ( .A1(n2972), .A2(n2687), .B1(n2971), .B2(n2970), .ZN(n2973)
         );
  INV_X4 U1305 ( .A(n2973), .ZN(n2980) );
  NAND2_X2 U1306 ( .A1(n3049), .A2(n2975), .ZN(n2974) );
  NAND2_X2 U1307 ( .A1(n3051), .A2(n2975), .ZN(n2976) );
  OAI221_X2 U1308 ( .B1(n454), .B2(n3055), .C1(n346), .C2(n3053), .A(n2976), 
        .ZN(n1267) );
  INV_X4 U1309 ( .A(U3_U3_DATA6_5), .ZN(n2977) );
  OAI22_X2 U1310 ( .A1(n3038), .A2(n2977), .B1(n283), .B2(n3036), .ZN(n1345)
         );
  INV_X4 U1311 ( .A(n2978), .ZN(n2981) );
  NOR2_X2 U1312 ( .A1(n2557), .A2(n2978), .ZN(n2979) );
  OAI22_X2 U1313 ( .A1(n2981), .A2(n2687), .B1(n2980), .B2(n2979), .ZN(n2982)
         );
  INV_X4 U1314 ( .A(n2982), .ZN(n2989) );
  NAND2_X2 U1315 ( .A1(n3049), .A2(n2984), .ZN(n2983) );
  NAND2_X2 U1316 ( .A1(n3051), .A2(n2984), .ZN(n2985) );
  OAI221_X2 U1317 ( .B1(n453), .B2(n3055), .C1(n345), .C2(n3053), .A(n2985), 
        .ZN(n1266) );
  INV_X4 U1318 ( .A(U3_U3_DATA6_6), .ZN(n2986) );
  OAI22_X2 U1319 ( .A1(n3038), .A2(n2986), .B1(n281), .B2(n3036), .ZN(n1344)
         );
  INV_X4 U1320 ( .A(n2987), .ZN(n2990) );
  NOR2_X2 U1321 ( .A1(n2557), .A2(n2987), .ZN(n2988) );
  OAI22_X2 U1322 ( .A1(n2990), .A2(n2687), .B1(n2989), .B2(n2988), .ZN(n2991)
         );
  INV_X4 U1323 ( .A(n2991), .ZN(n2998) );
  NAND2_X2 U1324 ( .A1(n3049), .A2(n2993), .ZN(n2992) );
  NAND2_X2 U1325 ( .A1(n3051), .A2(n2993), .ZN(n2994) );
  OAI221_X2 U1326 ( .B1(n452), .B2(n3055), .C1(n344), .C2(n3053), .A(n2994), 
        .ZN(n1265) );
  INV_X4 U1327 ( .A(U3_U3_DATA6_7), .ZN(n2995) );
  OAI22_X2 U1328 ( .A1(n3038), .A2(n2995), .B1(n279), .B2(n3036), .ZN(n1343)
         );
  INV_X4 U1329 ( .A(n2996), .ZN(n2999) );
  NOR2_X2 U1330 ( .A1(n2557), .A2(n2996), .ZN(n2997) );
  OAI22_X2 U1331 ( .A1(n2999), .A2(n2687), .B1(n2998), .B2(n2997), .ZN(n3000)
         );
  NAND2_X2 U1332 ( .A1(n3049), .A2(n3002), .ZN(n3001) );
  NAND2_X2 U1333 ( .A1(n3051), .A2(n3002), .ZN(n3003) );
  OAI221_X2 U1334 ( .B1(n451), .B2(n3055), .C1(n343), .C2(n3053), .A(n3003), 
        .ZN(n1264) );
  INV_X4 U1335 ( .A(U3_U3_DATA6_8), .ZN(n3004) );
  OAI22_X2 U1336 ( .A1(n3038), .A2(n3004), .B1(n277), .B2(n3036), .ZN(n1326)
         );
  NAND2_X2 U1337 ( .A1(n3049), .A2(n3007), .ZN(n3006) );
  NAND2_X2 U1338 ( .A1(n3051), .A2(n3007), .ZN(n3008) );
  OAI221_X2 U1339 ( .B1(n450), .B2(n3055), .C1(n342), .C2(n3053), .A(n3008), 
        .ZN(n1263) );
  INV_X4 U1340 ( .A(U3_U3_DATA6_9), .ZN(n3009) );
  OAI22_X2 U1341 ( .A1(n3038), .A2(n3009), .B1(n275), .B2(n3036), .ZN(n1325)
         );
  INV_X4 U1342 ( .A(n3010), .ZN(n3012) );
  NOR2_X2 U1343 ( .A1(n2557), .A2(n3010), .ZN(n3011) );
  OAI22_X2 U1344 ( .A1(n3012), .A2(n2687), .B1(n2604), .B2(n3011), .ZN(n3013)
         );
  INV_X4 U1345 ( .A(n3013), .ZN(n3020) );
  NAND2_X2 U1346 ( .A1(n3049), .A2(n3015), .ZN(n3014) );
  OAI221_X2 U1347 ( .B1(n275), .B2(net10950), .C1(n17), .C2(net10887), .A(
        n3014), .ZN(n1275) );
  NAND2_X2 U1348 ( .A1(n3051), .A2(n3015), .ZN(n3016) );
  OAI221_X2 U1349 ( .B1(n449), .B2(n3055), .C1(n341), .C2(n3053), .A(n3016), 
        .ZN(n1262) );
  INV_X4 U1350 ( .A(U3_U3_DATA6_10), .ZN(n3017) );
  OAI22_X2 U1351 ( .A1(n3038), .A2(n3017), .B1(n273), .B2(n3036), .ZN(n1324)
         );
  INV_X4 U1352 ( .A(n3018), .ZN(n3021) );
  NOR2_X2 U1353 ( .A1(n2557), .A2(n3018), .ZN(n3019) );
  OAI22_X2 U1354 ( .A1(n3021), .A2(n2687), .B1(n3020), .B2(n3019), .ZN(n3022)
         );
  INV_X4 U1355 ( .A(n3022), .ZN(n3029) );
  NAND2_X2 U1356 ( .A1(n3049), .A2(n3024), .ZN(n3023) );
  OAI221_X2 U1357 ( .B1(n273), .B2(net10950), .C1(n15), .C2(net10887), .A(
        n3023), .ZN(n1274) );
  NAND2_X2 U1358 ( .A1(n3051), .A2(n3024), .ZN(n3025) );
  OAI221_X2 U1359 ( .B1(n448), .B2(n3055), .C1(n340), .C2(n3053), .A(n3025), 
        .ZN(n1261) );
  XNOR2_X2 U1360 ( .A(r520_carry[11]), .B(graphRead1_Addr[11]), .ZN(n3026) );
  OAI22_X2 U1361 ( .A1(n3038), .A2(n3026), .B1(n271), .B2(n3036), .ZN(n1323)
         );
  INV_X4 U1362 ( .A(n3027), .ZN(n3030) );
  NOR2_X2 U1363 ( .A1(n2557), .A2(n3027), .ZN(n3028) );
  OAI22_X2 U1364 ( .A1(n3030), .A2(n2687), .B1(n3029), .B2(n3028), .ZN(n3031)
         );
  INV_X4 U1365 ( .A(n3031), .ZN(n3043) );
  NAND2_X2 U1366 ( .A1(n3049), .A2(n3033), .ZN(n3032) );
  OAI221_X2 U1367 ( .B1(n271), .B2(net10950), .C1(n13), .C2(net10887), .A(
        n3032), .ZN(n1273) );
  INV_X4 U1368 ( .A(graphRead1_DataInput[11]), .ZN(n3035) );
  NAND2_X2 U1369 ( .A1(n3051), .A2(n3033), .ZN(n3034) );
  OAI221_X2 U1370 ( .B1(n3055), .B2(n3035), .C1(n339), .C2(n3053), .A(n3034), 
        .ZN(n1260) );
  NAND2_X2 U1371 ( .A1(graphRead1_Addr[11]), .A2(r520_carry[11]), .ZN(n3037)
         );
  NOR2_X2 U1372 ( .A1(n3038), .A2(n3037), .ZN(n3039) );
  MUX2_X2 U1373 ( .A(n3040), .B(n3039), .S(n270), .Z(n1322) );
  INV_X4 U1374 ( .A(n3041), .ZN(n3044) );
  NOR2_X2 U1375 ( .A1(n2557), .A2(n3041), .ZN(n3042) );
  OAI22_X2 U1376 ( .A1(n3044), .A2(n2687), .B1(n3043), .B2(n3042), .ZN(n3048)
         );
  XOR2_X2 U1377 ( .A(n2687), .B(n3046), .Z(n3047) );
  NAND2_X2 U1378 ( .A1(n3049), .A2(n2657), .ZN(n3050) );
  OAI221_X2 U1379 ( .B1(n270), .B2(net10950), .C1(n11), .C2(net10887), .A(
        n3050), .ZN(n1272) );
  INV_X4 U1380 ( .A(graphRead1_DataInput[12]), .ZN(n3054) );
  NAND2_X2 U1381 ( .A1(n3051), .A2(n2657), .ZN(n3052) );
  OAI221_X2 U1382 ( .B1(n3055), .B2(n3054), .C1(n338), .C2(n3053), .A(n3052), 
        .ZN(n1259) );
  NAND2_X2 U1383 ( .A1(net10942), .A2(net10943), .ZN(n3116) );
  INV_X4 U1384 ( .A(n3116), .ZN(n3157) );
  XOR2_X2 U1385 ( .A(U3_U6_Z_0), .B(net10840), .Z(net10940) );
  INV_X4 U1386 ( .A(n267), .ZN(net10939) );
  NAND2_X2 U1387 ( .A1(n2573), .A2(net10939), .ZN(n3056) );
  OAI221_X2 U1388 ( .B1(n336), .B2(n3068), .C1(n473), .C2(n2565), .A(n3056), 
        .ZN(n1403) );
  XOR2_X2 U1389 ( .A(net10931), .B(net10840), .Z(n3057) );
  XOR2_X2 U1390 ( .A(n3057), .B(net10927), .Z(n265) );
  XOR2_X2 U1391 ( .A(net10923), .B(net10840), .Z(n3058) );
  XOR2_X2 U1392 ( .A(n3058), .B(net10919), .Z(n263) );
  XOR2_X2 U1393 ( .A(net10915), .B(net10840), .Z(n3059) );
  XOR2_X2 U1394 ( .A(n3059), .B(net10911), .Z(n261) );
  XOR2_X2 U1395 ( .A(net10907), .B(net10840), .Z(n3060) );
  XOR2_X2 U1396 ( .A(n3060), .B(net10903), .Z(n259) );
  INV_X4 U1397 ( .A(n259), .ZN(n3061) );
  NAND2_X2 U1398 ( .A1(n2573), .A2(n3061), .ZN(n3062) );
  OAI221_X2 U1399 ( .B1(n332), .B2(n3068), .C1(n469), .C2(n2565), .A(n3062), 
        .ZN(n1399) );
  XOR2_X2 U1400 ( .A(net10899), .B(net10840), .Z(n3063) );
  INV_X4 U1401 ( .A(n257), .ZN(n3064) );
  NAND2_X2 U1402 ( .A1(n2573), .A2(n3064), .ZN(n3065) );
  OAI221_X2 U1403 ( .B1(n331), .B2(n3068), .C1(n468), .C2(n2565), .A(n3065), 
        .ZN(n1398) );
  XOR2_X2 U1404 ( .A(net10893), .B(net10844), .Z(n255) );
  INV_X4 U1405 ( .A(n255), .ZN(n3066) );
  NAND2_X2 U1406 ( .A1(n2573), .A2(n3066), .ZN(n3067) );
  OAI221_X2 U1407 ( .B1(n294), .B2(n3068), .C1(n467), .C2(n2565), .A(n3067), 
        .ZN(n1397) );
  INV_X4 U1408 ( .A(net10887), .ZN(net10885) );
  NAND2_X2 U1409 ( .A1(net10884), .A2(net10867), .ZN(n3071) );
  OAI221_X2 U1410 ( .B1(net10881), .B2(n293), .C1(n87), .C2(n3084), .A(n3070), 
        .ZN(n1334) );
  INV_X4 U1411 ( .A(net10881), .ZN(net10863) );
  INV_X4 U1412 ( .A(n3071), .ZN(n3086) );
  INV_X4 U1413 ( .A(n3073), .ZN(n1333) );
  INV_X4 U1414 ( .A(n3075), .ZN(n1332) );
  INV_X4 U1415 ( .A(n3077), .ZN(n1328) );
  INV_X4 U1416 ( .A(n3079), .ZN(n1327) );
  INV_X4 U1417 ( .A(n3081), .ZN(n1329) );
  INV_X4 U1418 ( .A(n3083), .ZN(n1330) );
  INV_X4 U1419 ( .A(n3087), .ZN(n1331) );
  NAND4_X2 U1420 ( .A1(n15), .A2(n31), .A3(n11), .A4(n13), .ZN(n1067) );
  INV_X4 U1421 ( .A(inputSRAM_Data[0]), .ZN(n3090) );
  INV_X4 U1422 ( .A(inputSRAM_Data[1]), .ZN(n3089) );
  INV_X4 U1423 ( .A(inputSRAM_Data[2]), .ZN(n3088) );
  INV_X4 U1424 ( .A(n424), .ZN(n3091) );
  NAND2_X2 U1425 ( .A1(n2581), .A2(n3093), .ZN(n3094) );
  NAND2_X2 U1426 ( .A1(reset), .A2(n3094), .ZN(n1051) );
  XNOR2_X2 U1427 ( .A(net10840), .B(net10839), .ZN(net10842) );
  INV_X4 U1428 ( .A(n3095), .ZN(n3097) );
  NAND3_X2 U1429 ( .A1(n3097), .A2(n3113), .A3(n845), .ZN(n54) );
  INV_X4 U1430 ( .A(n54), .ZN(n991) );
  NOR2_X2 U1431 ( .A1(n3113), .A2(n3098), .ZN(n3099) );
  AOI221_X2 U1432 ( .B1(U97_DATA2_0), .B2(n3115), .C1(U97_DATA4_0), .C2(n564), 
        .A(n3099), .ZN(n1005) );
  NOR2_X2 U1433 ( .A1(n3113), .A2(n3100), .ZN(n3101) );
  AOI221_X2 U1434 ( .B1(U97_DATA2_1), .B2(n3115), .C1(U97_DATA4_1), .C2(n564), 
        .A(n3101), .ZN(n1003) );
  NOR2_X2 U1435 ( .A1(n3113), .A2(n3102), .ZN(n3103) );
  AOI221_X2 U1436 ( .B1(U97_DATA2_2), .B2(n3115), .C1(U97_DATA4_2), .C2(n564), 
        .A(n3103), .ZN(n1001) );
  NOR2_X2 U1437 ( .A1(n3113), .A2(n3104), .ZN(n3105) );
  AOI221_X2 U1438 ( .B1(U97_DATA2_3), .B2(n3115), .C1(U97_DATA4_3), .C2(n564), 
        .A(n3105), .ZN(n999) );
  NOR2_X2 U1439 ( .A1(n3113), .A2(n3106), .ZN(n3107) );
  AOI221_X2 U1440 ( .B1(U97_DATA2_4), .B2(n3115), .C1(U97_DATA4_4), .C2(n564), 
        .A(n3107), .ZN(n997) );
  NOR2_X2 U1441 ( .A1(n3113), .A2(n3108), .ZN(n3109) );
  AOI221_X2 U1442 ( .B1(U97_DATA2_5), .B2(n3115), .C1(U97_DATA4_5), .C2(n564), 
        .A(n3109), .ZN(n995) );
  NOR2_X2 U1443 ( .A1(n3113), .A2(n3110), .ZN(n3111) );
  AOI221_X2 U1444 ( .B1(U97_DATA2_6), .B2(n3115), .C1(U97_DATA4_6), .C2(n564), 
        .A(n3111), .ZN(n993) );
  NOR2_X2 U1445 ( .A1(n3113), .A2(n3112), .ZN(n3114) );
  AOI221_X2 U1446 ( .B1(U97_DATA2_7), .B2(n3115), .C1(U97_DATA4_7), .C2(n564), 
        .A(n3114), .ZN(n988) );
  INV_X4 U1447 ( .A(n831), .ZN(n70) );
  OAI22_X2 U1448 ( .A1(n506), .A2(net11668), .B1(n178), .B2(net11700), .ZN(
        n1240) );
  OAI22_X2 U1449 ( .A1(n490), .A2(net11668), .B1(n162), .B2(net11694), .ZN(
        n1256) );
  OAI22_X2 U1450 ( .A1(n482), .A2(net11668), .B1(n146), .B2(net11700), .ZN(
        n1168) );
  OAI22_X2 U1451 ( .A1(n466), .A2(net11670), .B1(n111), .B2(net11696), .ZN(
        n1176) );
  OAI22_X2 U1452 ( .A1(n538), .A2(net11668), .B1(n226), .B2(net11696), .ZN(
        n1208) );
  OAI22_X2 U1453 ( .A1(n554), .A2(net11670), .B1(n242), .B2(net11696), .ZN(
        n1192) );
  OAI22_X2 U1454 ( .A1(n522), .A2(net11670), .B1(n194), .B2(net11696), .ZN(
        n1224) );
  OAI22_X2 U1455 ( .A1(n530), .A2(net11668), .B1(n210), .B2(net11696), .ZN(
        n1216) );
  OAI22_X2 U1456 ( .A1(n505), .A2(net11670), .B1(n177), .B2(net11696), .ZN(
        n1241) );
  OAI22_X2 U1457 ( .A1(n489), .A2(net11668), .B1(n161), .B2(net11696), .ZN(
        n1257) );
  OAI22_X2 U1458 ( .A1(n481), .A2(net11668), .B1(n145), .B2(net11696), .ZN(
        n1169) );
  OAI22_X2 U1459 ( .A1(n465), .A2(net11670), .B1(n110), .B2(net11696), .ZN(
        n1177) );
  OAI22_X2 U1460 ( .A1(n537), .A2(net11670), .B1(n225), .B2(net11696), .ZN(
        n1209) );
  OAI22_X2 U1461 ( .A1(n553), .A2(net11668), .B1(n241), .B2(net11696), .ZN(
        n1193) );
  OAI22_X2 U1462 ( .A1(n521), .A2(net11668), .B1(n193), .B2(net11696), .ZN(
        n1225) );
  OAI22_X2 U1463 ( .A1(n529), .A2(net11668), .B1(n209), .B2(net11694), .ZN(
        n1217) );
  OAI22_X2 U1464 ( .A1(n504), .A2(net11670), .B1(n176), .B2(net11700), .ZN(
        n1242) );
  OAI22_X2 U1466 ( .A1(n480), .A2(net11670), .B1(n144), .B2(net11694), .ZN(
        n1170) );
  OAI22_X2 U1468 ( .A1(n536), .A2(net11670), .B1(n224), .B2(net11700), .ZN(
        n1210) );
  OAI22_X2 U1469 ( .A1(n552), .A2(net11668), .B1(n240), .B2(net11700), .ZN(
        n1194) );
  OAI22_X2 U1472 ( .A1(n503), .A2(net11668), .B1(n175), .B2(net11700), .ZN(
        n1243) );
  OAI22_X2 U1474 ( .A1(n479), .A2(net11670), .B1(n143), .B2(net11694), .ZN(
        n1171) );
  OAI22_X2 U1475 ( .A1(n463), .A2(net11670), .B1(n108), .B2(net11694), .ZN(
        n1179) );
  OAI22_X2 U1476 ( .A1(n535), .A2(net11668), .B1(n223), .B2(net11700), .ZN(
        n1211) );
  OAI22_X2 U1477 ( .A1(n551), .A2(net11670), .B1(n239), .B2(net11694), .ZN(
        n1195) );
  OAI22_X2 U1478 ( .A1(n519), .A2(net11668), .B1(n191), .B2(net11700), .ZN(
        n1227) );
  OAI22_X2 U1479 ( .A1(n527), .A2(net11668), .B1(n207), .B2(net11694), .ZN(
        n1219) );
  OAI22_X2 U1480 ( .A1(n502), .A2(net11670), .B1(n174), .B2(net11700), .ZN(
        n1244) );
  OAI22_X2 U1481 ( .A1(n486), .A2(net10805), .B1(n158), .B2(net11694), .ZN(
        n1164) );
  OAI22_X2 U1482 ( .A1(n478), .A2(net11670), .B1(n142), .B2(net11700), .ZN(
        n1172) );
  OAI22_X2 U1483 ( .A1(n462), .A2(net11668), .B1(n107), .B2(net11694), .ZN(
        n1180) );
  OAI22_X2 U1484 ( .A1(n534), .A2(net11670), .B1(n222), .B2(net11700), .ZN(
        n1212) );
  OAI22_X2 U1485 ( .A1(n550), .A2(net11668), .B1(n238), .B2(net11694), .ZN(
        n1196) );
  OAI22_X2 U1486 ( .A1(n518), .A2(net11668), .B1(n190), .B2(net11700), .ZN(
        n1228) );
  OAI22_X2 U1487 ( .A1(n526), .A2(net10805), .B1(n206), .B2(net11700), .ZN(
        n1220) );
  OAI22_X2 U1488 ( .A1(n501), .A2(net10805), .B1(n173), .B2(net11694), .ZN(
        n1245) );
  OAI22_X2 U1489 ( .A1(n485), .A2(net11670), .B1(n157), .B2(net11700), .ZN(
        n1165) );
  OAI22_X2 U1490 ( .A1(n477), .A2(net11668), .B1(n141), .B2(net11694), .ZN(
        n1173) );
  OAI22_X2 U1491 ( .A1(n461), .A2(net10805), .B1(n106), .B2(net11700), .ZN(
        n1181) );
  OAI22_X2 U1492 ( .A1(n533), .A2(net11668), .B1(n221), .B2(net11694), .ZN(
        n1213) );
  OAI22_X2 U1493 ( .A1(n549), .A2(net11670), .B1(n237), .B2(net11700), .ZN(
        n1197) );
  OAI22_X2 U1494 ( .A1(n517), .A2(net10805), .B1(n189), .B2(net11694), .ZN(
        n1229) );
  OAI22_X2 U1495 ( .A1(n525), .A2(net10805), .B1(n205), .B2(net11700), .ZN(
        n1221) );
  OAI22_X2 U1496 ( .A1(n500), .A2(net10805), .B1(n172), .B2(net11694), .ZN(
        n1246) );
  OAI22_X2 U1497 ( .A1(n484), .A2(net11670), .B1(n156), .B2(net11700), .ZN(
        n1166) );
  OAI22_X2 U1498 ( .A1(n476), .A2(net11668), .B1(n140), .B2(net11694), .ZN(
        n1174) );
  OAI22_X2 U1499 ( .A1(n460), .A2(net10805), .B1(n105), .B2(net11700), .ZN(
        n1182) );
  OAI22_X2 U1500 ( .A1(n532), .A2(net10805), .B1(n220), .B2(net11694), .ZN(
        n1214) );
  OAI22_X2 U1501 ( .A1(n548), .A2(net11670), .B1(n236), .B2(net11696), .ZN(
        n1198) );
  OAI22_X2 U1502 ( .A1(n516), .A2(net10805), .B1(n188), .B2(net11694), .ZN(
        n1230) );
  OAI22_X2 U1503 ( .A1(n524), .A2(net11670), .B1(n204), .B2(net11696), .ZN(
        n1222) );
  OAI22_X2 U1504 ( .A1(n499), .A2(net10805), .B1(n171), .B2(net11700), .ZN(
        n1247) );
  OAI22_X2 U1505 ( .A1(n483), .A2(net11670), .B1(n155), .B2(net11694), .ZN(
        n1167) );
  OAI22_X2 U1506 ( .A1(n475), .A2(net11670), .B1(n139), .B2(net11700), .ZN(
        n1175) );
  OAI22_X2 U1507 ( .A1(n459), .A2(net10805), .B1(n104), .B2(net11694), .ZN(
        n1183) );
  OAI22_X2 U1508 ( .A1(n531), .A2(net10805), .B1(n219), .B2(net11700), .ZN(
        n1215) );
  OAI22_X2 U1509 ( .A1(n547), .A2(net10805), .B1(n235), .B2(net11700), .ZN(
        n1199) );
  OAI22_X2 U1510 ( .A1(n515), .A2(net10805), .B1(n187), .B2(net11694), .ZN(
        n1231) );
  OAI22_X2 U1511 ( .A1(n523), .A2(net11668), .B1(n203), .B2(net11696), .ZN(
        n1223) );
  AOI221_X2 U1512 ( .B1(U38_DATA5_0), .B2(n2471), .C1(U38_DATA6_0), .C2(n2472), 
        .A(n3117), .ZN(n3120) );
  NAND2_X2 U1513 ( .A1(n3120), .A2(n3119), .ZN(n3121) );
  NAND2_X2 U1514 ( .A1(n2653), .A2(n3121), .ZN(n630) );
  AOI221_X2 U1515 ( .B1(U38_DATA5_1), .B2(n2471), .C1(U38_DATA6_1), .C2(n2472), 
        .A(n3122), .ZN(n3125) );
  NAND2_X2 U1516 ( .A1(n3125), .A2(n3124), .ZN(n3126) );
  NAND2_X2 U1517 ( .A1(n2653), .A2(n3126), .ZN(n624) );
  AOI221_X2 U1518 ( .B1(U38_DATA5_2), .B2(n2471), .C1(U38_DATA6_2), .C2(n2472), 
        .A(n3127), .ZN(n3130) );
  NAND2_X2 U1519 ( .A1(n3130), .A2(n3129), .ZN(n3131) );
  NAND2_X2 U1520 ( .A1(n2653), .A2(n3131), .ZN(n618) );
  AOI221_X2 U1521 ( .B1(U38_DATA5_3), .B2(n2471), .C1(U38_DATA6_3), .C2(n2472), 
        .A(n3132), .ZN(n3135) );
  NAND2_X2 U1522 ( .A1(n3135), .A2(n3134), .ZN(n3136) );
  NAND2_X2 U1523 ( .A1(n2653), .A2(n3136), .ZN(n612) );
  AOI221_X2 U1524 ( .B1(U38_DATA5_4), .B2(n2471), .C1(U38_DATA6_4), .C2(n2472), 
        .A(n3137), .ZN(n3140) );
  NAND2_X2 U1525 ( .A1(n3140), .A2(n3139), .ZN(n3141) );
  NAND2_X2 U1526 ( .A1(n2653), .A2(n3141), .ZN(n606) );
  AOI221_X2 U1527 ( .B1(U38_DATA5_5), .B2(n2471), .C1(U38_DATA6_5), .C2(n2472), 
        .A(n3142), .ZN(n3145) );
  NAND2_X2 U1528 ( .A1(n3145), .A2(n3144), .ZN(n3146) );
  NAND2_X2 U1529 ( .A1(n2653), .A2(n3146), .ZN(n600) );
  AOI221_X2 U1530 ( .B1(U38_DATA5_6), .B2(n2471), .C1(U38_DATA6_6), .C2(n2472), 
        .A(n3147), .ZN(n3150) );
  NAND2_X2 U1531 ( .A1(n3150), .A2(n3149), .ZN(n3151) );
  NAND2_X2 U1532 ( .A1(n2653), .A2(n3151), .ZN(n594) );
  AOI221_X2 U1533 ( .B1(U38_DATA5_7), .B2(n2471), .C1(U38_DATA6_7), .C2(n2472), 
        .A(n3152), .ZN(n3155) );
  NAND2_X2 U1534 ( .A1(n3155), .A2(n3154), .ZN(n3156) );
  NAND2_X2 U1535 ( .A1(n2653), .A2(n3156), .ZN(n578) );
  NAND2_X2 U3 ( .A1(n682), .A2(reset), .ZN(n1047) );
  NAND2_X2 U4 ( .A1(n2687), .A2(net11093), .ZN(net10887) );
  OAI22_X1 U5 ( .A1(n488), .A2(net10805), .B1(n160), .B2(net11700), .ZN(n1258)
         );
  OAI22_X1 U6 ( .A1(n464), .A2(net10805), .B1(n109), .B2(net11694), .ZN(n1178)
         );
  OAI22_X1 U7 ( .A1(n520), .A2(net10805), .B1(n192), .B2(net11694), .ZN(n1226)
         );
  OAI22_X1 U8 ( .A1(n528), .A2(net10805), .B1(n208), .B2(net11694), .ZN(n1218)
         );
  OAI22_X1 U9 ( .A1(n487), .A2(net10805), .B1(n159), .B2(net11700), .ZN(n1163)
         );
  INV_X8 U10 ( .A(net11682), .ZN(net11668) );
  INV_X8 U11 ( .A(net11682), .ZN(net11670) );
endmodule


module fsm ( clock, reset, start, graphData1_Zero, iterDone, iterStop, 
        negCycle, zeroFlag, outputWriteDone, goS8, fsm_state );
  output [4:0] fsm_state;
  input clock, reset, start, graphData1_Zero, iterDone, iterStop, negCycle,
         zeroFlag, outputWriteDone, goS8;
  wire   U9_Z_0, U9_Z_3, U9_Z_4, n15, n16, n18, n23, n55, net10661, net10662,
         net10663, net10665, net10670, net10678, net10680, net10682, net10683,
         net10685, net10690, net10693, net10707, net10709, net10714, net10715,
         net10719, net10720, net10721, net10722, net10739, net10744, net10745,
         net10746, net12553, net12554, net12555, net17856, net17866, net10718,
         net12636, net12552, net10692, n222, n223, n224, n225, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264;
  wire   [175:171] n;

  INV_X4 U76 ( .A(negCycle), .ZN(n23) );
  DFF_X2 current_state_reg_4_ ( .D(U9_Z_4), .CK(clock), .Q(n[175]), .QN(
        net10739) );
  DFF_X2 current_state_reg_0_ ( .D(U9_Z_0), .CK(clock), .Q(n[171]), .QN(n18)
         );
  SDFF_X1 current_state_reg_2_ ( .D(reset), .SI(1'b0), .SE(n55), .CK(clock), 
        .Q(n[173]), .QN(n16) );
  DFF_X2 current_state_reg_3_ ( .D(U9_Z_3), .CK(clock), .Q(n[174]), .QN(n15)
         );
  SDFF_X2 current_state_reg_1_ ( .D(reset), .SI(1'b0), .SE(n238), .CK(clock), 
        .Q(n[172]), .QN(net10746) );
  NAND4_X2 U3 ( .A1(n264), .A2(n240), .A3(n243), .A4(n244), .ZN(fsm_state[4])
         );
  NOR2_X2 U4 ( .A1(n[174]), .A2(n18), .ZN(net12555) );
  NOR2_X2 U5 ( .A1(n18), .A2(n15), .ZN(net17856) );
  OAI211_X2 U6 ( .C1(n222), .C2(net10692), .A(net10720), .B(n243), .ZN(n252)
         );
  INV_X4 U7 ( .A(net12555), .ZN(n222) );
  NOR2_X2 U8 ( .A1(n15), .A2(net10692), .ZN(net12636) );
  OR3_X4 U9 ( .A1(net10661), .A2(negCycle), .A3(iterStop), .ZN(n233) );
  OAI211_X2 U10 ( .C1(n250), .C2(net10709), .A(n240), .B(net10721), .ZN(n223)
         );
  INV_X4 U11 ( .A(n223), .ZN(n241) );
  NAND4_X1 U12 ( .A1(n235), .A2(n[173]), .A3(net10746), .A4(n[175]), .ZN(n240)
         );
  NAND3_X1 U13 ( .A1(n225), .A2(net10665), .A3(net10715), .ZN(net10714) );
  OR2_X4 U14 ( .A1(n264), .A2(zeroFlag), .ZN(n245) );
  AOI21_X2 U15 ( .B1(start), .B2(n224), .A(net10690), .ZN(n251) );
  INV_X4 U16 ( .A(net10692), .ZN(n224) );
  OAI21_X2 U17 ( .B1(negCycle), .B2(iterStop), .A(net10678), .ZN(net10715) );
  NOR3_X2 U18 ( .A1(n16), .A2(n[175]), .A3(net10746), .ZN(net12554) );
  OAI33_X1 U19 ( .A1(n[174]), .A2(n[171]), .A3(n251), .B1(net10661), .B2(
        iterStop), .B3(n23), .ZN(net10683) );
  NAND4_X2 U20 ( .A1(n257), .A2(n259), .A3(n256), .A4(net10663), .ZN(
        fsm_state[0]) );
  NAND3_X1 U21 ( .A1(n16), .A2(net10746), .A3(net10739), .ZN(net10692) );
  AND2_X4 U22 ( .A1(net12636), .A2(n18), .ZN(net12552) );
  NOR2_X2 U23 ( .A1(net10722), .A2(net12552), .ZN(net10718) );
  NOR4_X2 U24 ( .A1(net10682), .A2(net10683), .A3(net12552), .A4(net10685), 
        .ZN(net10680) );
  NAND2_X2 U25 ( .A1(net12636), .A2(n[171]), .ZN(net10720) );
  NAND4_X2 U26 ( .A1(n225), .A2(net10661), .A3(net10662), .A4(net10663), .ZN(
        fsm_state[3]) );
  AND4_X2 U27 ( .A1(net10718), .A2(net10719), .A3(net10720), .A4(net10721), 
        .ZN(n225) );
  NAND2_X2 U28 ( .A1(net17866), .A2(net17856), .ZN(net10661) );
  NAND2_X2 U29 ( .A1(net12554), .A2(net17856), .ZN(net10662) );
  NAND2_X2 U30 ( .A1(net10690), .A2(net17856), .ZN(net10663) );
  INV_X4 U31 ( .A(net10670), .ZN(net10722) );
  NAND2_X2 U32 ( .A1(net12554), .A2(net12553), .ZN(net10719) );
  NAND2_X2 U33 ( .A1(net10690), .A2(net12553), .ZN(net10721) );
  NOR3_X2 U34 ( .A1(n228), .A2(n253), .A3(net10678), .ZN(n254) );
  NOR4_X1 U35 ( .A1(n237), .A2(net10707), .A3(n252), .A4(net10685), .ZN(n238)
         );
  NAND2_X1 U36 ( .A1(n229), .A2(n[172]), .ZN(n258) );
  NOR4_X1 U37 ( .A1(n228), .A2(n230), .A3(net10678), .A4(n261), .ZN(n55) );
  AND3_X4 U38 ( .A1(n16), .A2(net10739), .A3(n[172]), .ZN(net17866) );
  NAND2_X1 U41 ( .A1(n260), .A2(n236), .ZN(net10685) );
  NAND3_X1 U42 ( .A1(net10746), .A2(n[171]), .A3(n229), .ZN(n243) );
  AND2_X4 U43 ( .A1(n[174]), .A2(n18), .ZN(net12553) );
  AOI21_X1 U44 ( .B1(net17866), .B2(n235), .A(n239), .ZN(n260) );
  AND2_X1 U45 ( .A1(net12555), .A2(net17866), .ZN(n228) );
  INV_X4 U46 ( .A(reset), .ZN(n231) );
  NOR3_X2 U47 ( .A1(n[174]), .A2(net10739), .A3(n[173]), .ZN(n229) );
  AND2_X1 U48 ( .A1(zeroFlag), .A2(n253), .ZN(n230) );
  INV_X4 U49 ( .A(net10662), .ZN(net10744) );
  NAND3_X2 U50 ( .A1(n[172]), .A2(n[171]), .A3(n229), .ZN(n264) );
  INV_X4 U51 ( .A(n264), .ZN(n253) );
  NAND3_X2 U52 ( .A1(net10739), .A2(net10746), .A3(n[173]), .ZN(net10709) );
  INV_X4 U53 ( .A(net10709), .ZN(net10690) );
  INV_X4 U54 ( .A(net10663), .ZN(net10745) );
  NAND2_X2 U55 ( .A1(n15), .A2(n18), .ZN(n250) );
  INV_X4 U56 ( .A(n250), .ZN(n235) );
  NAND2_X2 U57 ( .A1(n18), .A2(n229), .ZN(n244) );
  NAND3_X2 U58 ( .A1(n240), .A2(n243), .A3(n244), .ZN(n263) );
  NOR4_X2 U59 ( .A1(net10744), .A2(n230), .A3(net10745), .A4(n263), .ZN(n232)
         );
  NOR2_X2 U60 ( .A1(n232), .A2(n231), .ZN(U9_Z_4) );
  NAND2_X2 U61 ( .A1(net12553), .A2(net17866), .ZN(net10670) );
  NAND2_X2 U62 ( .A1(net12555), .A2(net10690), .ZN(n256) );
  INV_X4 U63 ( .A(graphData1_Zero), .ZN(n247) );
  INV_X4 U64 ( .A(net10661), .ZN(net10678) );
  OAI221_X2 U65 ( .B1(goS8), .B2(net10670), .C1(n256), .C2(n247), .A(n233), 
        .ZN(n237) );
  INV_X4 U66 ( .A(net10721), .ZN(net10707) );
  NAND2_X2 U67 ( .A1(net12554), .A2(n235), .ZN(n234) );
  NAND2_X2 U68 ( .A1(n234), .A2(net10719), .ZN(n239) );
  NAND2_X2 U69 ( .A1(iterDone), .A2(net10722), .ZN(n236) );
  NAND2_X2 U70 ( .A1(net12555), .A2(net12554), .ZN(net10665) );
  AND2_X1 U71 ( .A1(reset), .A2(net10714), .ZN(U9_Z_3) );
  INV_X4 U72 ( .A(n239), .ZN(n242) );
  NAND4_X2 U73 ( .A1(n242), .A2(n256), .A3(net10663), .A4(n241), .ZN(n261) );
  INV_X4 U74 ( .A(n243), .ZN(n249) );
  INV_X4 U75 ( .A(n256), .ZN(n248) );
  NAND2_X2 U77 ( .A1(n245), .A2(n244), .ZN(n246) );
  AOI221_X2 U78 ( .B1(outputWriteDone), .B2(n249), .C1(n248), .C2(n247), .A(
        n246), .ZN(net10693) );
  INV_X4 U79 ( .A(net10693), .ZN(net10682) );
  NOR2_X2 U80 ( .A1(net10680), .A2(n231), .ZN(U9_Z_0) );
  INV_X4 U81 ( .A(n252), .ZN(n257) );
  NAND3_X2 U82 ( .A1(net10665), .A2(net10662), .A3(n254), .ZN(n255) );
  INV_X4 U83 ( .A(n255), .ZN(n259) );
  NAND4_X2 U84 ( .A1(n260), .A2(n259), .A3(n258), .A4(net10670), .ZN(
        fsm_state[1]) );
  INV_X4 U85 ( .A(n261), .ZN(n262) );
  NAND3_X2 U86 ( .A1(n262), .A2(net10665), .A3(net10662), .ZN(fsm_state[2]) );
endmodule


module top_without_mem ( clock, reset, start, inputSRAM_Data, 
        graphRead1_DataInput, graphRead2_DataInput, workRead1_DataInput, 
        workRead2_DataInput, inputSRAM_Addr, graphRead1_Addr, graphRead2_Addr, 
        workWrite_Dist, workWrite_Pred, workRead1_Addr, workRead2_Addr, 
        workWrite_Addr, work_WE, outputWrite_Data, outputWrite_Addr, output_WE
 );
  input [7:0] inputSRAM_Data;
  input [127:0] graphRead1_DataInput;
  input [127:0] graphRead2_DataInput;
  input [127:0] workRead1_DataInput;
  input [127:0] workRead2_DataInput;
  output [9:0] inputSRAM_Addr;
  output [12:0] graphRead1_Addr;
  output [12:0] graphRead2_Addr;
  output [16:0] workWrite_Dist;
  output [7:0] workWrite_Pred;
  output [12:0] workRead1_Addr;
  output [12:0] workRead2_Addr;
  output [12:0] workWrite_Addr;
  output [15:0] outputWrite_Data;
  output [13:0] outputWrite_Addr;
  input clock, reset, start;
  output work_WE, output_WE;
  wire   graphData1_Zero_reg, iterDone, iterStop, negCycle, zeroFlag,
         outputWriteDone, goS8, n32, n33, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15;
  wire   [4:0] state;

  datapath data ( .clock(clock), .reset(n32), .inputSRAM_Data(inputSRAM_Data), 
        .graphRead1_DataInput(graphRead1_DataInput), .graphRead2_DataInput(
        graphRead2_DataInput), .workRead1_DataInput(workRead1_DataInput), 
        .workRead2_DataInput(workRead2_DataInput), .inputSRAM_Addr(
        inputSRAM_Addr), .graphRead1_Addr(graphRead1_Addr), .graphRead2_Addr(
        graphRead2_Addr), .workWrite_Dist(workWrite_Dist), .workWrite_Pred(
        workWrite_Pred), .workRead1_Addr({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, 
        SYNOPSYS_UNCONNECTED_5, workRead1_Addr[7:0]}), .workRead2_Addr({
        SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, 
        SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, workRead2_Addr[7:0]}), 
        .workWrite_Addr({SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, 
        SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, 
        SYNOPSYS_UNCONNECTED_15, workWrite_Addr[7:0]}), .work_WE(work_WE), 
        .outputWrite_Data(outputWrite_Data), .outputWrite_Addr(
        outputWrite_Addr), .output_WE(output_WE), .state(state), 
        .graphData1_Zero_reg(graphData1_Zero_reg), .iterDone(iterDone), 
        .iterStop(iterStop), .negCycle(negCycle), .zeroFlag(zeroFlag), 
        .outputWriteDone(outputWriteDone), .goS8(goS8) );
  fsm control ( .clock(clock), .reset(n32), .start(start), .graphData1_Zero(
        graphData1_Zero_reg), .iterDone(iterDone), .iterStop(iterStop), 
        .negCycle(negCycle), .zeroFlag(zeroFlag), .outputWriteDone(
        outputWriteDone), .goS8(goS8), .fsm_state(state) );
  INV_X4 U1 ( .A(1'b1), .ZN(workWrite_Addr[8]) );
  INV_X4 U3 ( .A(1'b1), .ZN(workWrite_Addr[9]) );
  INV_X4 U5 ( .A(1'b1), .ZN(workWrite_Addr[10]) );
  INV_X4 U7 ( .A(1'b1), .ZN(workWrite_Addr[11]) );
  INV_X4 U9 ( .A(1'b1), .ZN(workWrite_Addr[12]) );
  INV_X4 U11 ( .A(1'b1), .ZN(workRead2_Addr[8]) );
  INV_X4 U13 ( .A(1'b1), .ZN(workRead2_Addr[9]) );
  INV_X4 U15 ( .A(1'b1), .ZN(workRead2_Addr[10]) );
  INV_X4 U17 ( .A(1'b1), .ZN(workRead2_Addr[11]) );
  INV_X4 U19 ( .A(1'b1), .ZN(workRead2_Addr[12]) );
  INV_X4 U21 ( .A(1'b1), .ZN(workRead1_Addr[8]) );
  INV_X4 U23 ( .A(1'b1), .ZN(workRead1_Addr[9]) );
  INV_X4 U25 ( .A(1'b1), .ZN(workRead1_Addr[10]) );
  INV_X4 U27 ( .A(1'b1), .ZN(workRead1_Addr[11]) );
  INV_X4 U29 ( .A(1'b1), .ZN(workRead1_Addr[12]) );
  INV_X4 U31 ( .A(n33), .ZN(n32) );
  INV_X4 U32 ( .A(reset), .ZN(n33) );
endmodule

